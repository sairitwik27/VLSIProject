magic
tech scmos
timestamp 1608917338
<< ab >>
rect 9 141 57 149
rect 18 76 57 141
rect 59 76 95 149
rect 18 13 55 76
rect 9 5 55 13
rect 57 5 95 76
rect 97 141 102 149
rect 97 85 99 141
rect 97 76 102 85
rect 104 76 167 149
rect 169 117 207 149
rect 169 76 216 117
rect 97 5 137 76
rect 139 5 202 76
rect 207 37 216 76
<< nwell >>
rect 0 37 216 117
<< pwell >>
rect 0 117 216 154
rect 0 0 216 37
<< poly >>
rect 26 136 28 141
rect 33 136 35 141
rect 46 134 48 138
rect 66 136 68 141
rect 73 136 75 141
rect 131 145 156 147
rect 114 140 116 145
rect 121 140 123 145
rect 86 134 88 138
rect 131 137 133 145
rect 141 137 143 141
rect 154 137 156 145
rect 154 135 159 137
rect 178 136 180 141
rect 185 136 187 141
rect 157 132 159 135
rect 26 112 28 125
rect 33 120 35 125
rect 46 120 48 125
rect 32 118 38 120
rect 32 116 34 118
rect 36 116 38 118
rect 32 114 38 116
rect 42 118 48 120
rect 42 116 44 118
rect 46 116 48 118
rect 42 114 48 116
rect 22 110 28 112
rect 22 108 24 110
rect 26 108 28 110
rect 22 106 28 108
rect 26 103 28 106
rect 36 103 38 114
rect 46 110 48 114
rect 66 112 68 125
rect 73 120 75 125
rect 86 120 88 125
rect 72 118 78 120
rect 72 116 74 118
rect 76 116 78 118
rect 72 114 78 116
rect 82 118 88 120
rect 114 119 116 128
rect 121 125 123 128
rect 121 123 125 125
rect 131 124 133 128
rect 141 125 143 128
rect 123 120 125 123
rect 141 123 150 125
rect 198 134 200 138
rect 141 121 146 123
rect 148 121 150 123
rect 82 116 84 118
rect 86 116 88 118
rect 82 114 88 116
rect 62 110 68 112
rect 62 108 64 110
rect 66 108 68 110
rect 62 106 68 108
rect 66 103 68 106
rect 76 103 78 114
rect 86 110 88 114
rect 113 117 119 119
rect 113 115 115 117
rect 117 115 119 117
rect 113 113 119 115
rect 123 118 129 120
rect 123 116 125 118
rect 127 116 129 118
rect 123 114 129 116
rect 141 119 150 121
rect 141 115 143 119
rect 157 115 159 123
rect 113 110 115 113
rect 123 110 125 114
rect 133 113 143 115
rect 149 113 162 115
rect 133 110 135 113
rect 149 110 151 113
rect 160 112 162 113
rect 178 112 180 125
rect 185 120 187 125
rect 198 120 200 125
rect 184 118 190 120
rect 184 116 186 118
rect 188 116 190 118
rect 184 114 190 116
rect 194 118 200 120
rect 194 116 196 118
rect 198 116 200 118
rect 194 114 200 116
rect 160 110 166 112
rect 26 85 28 90
rect 36 85 38 90
rect 46 88 48 92
rect 66 85 68 90
rect 76 85 78 90
rect 86 88 88 92
rect 123 88 125 92
rect 133 88 135 92
rect 113 79 115 83
rect 160 108 162 110
rect 164 108 166 110
rect 160 106 166 108
rect 174 110 180 112
rect 174 108 176 110
rect 178 108 180 110
rect 174 106 180 108
rect 178 103 180 106
rect 188 103 190 114
rect 198 110 200 114
rect 178 85 180 90
rect 188 85 190 90
rect 198 88 200 92
rect 149 79 151 83
rect 26 62 28 66
rect 36 64 38 69
rect 46 64 48 69
rect 66 64 68 69
rect 76 64 78 69
rect 155 71 157 75
rect 86 62 88 66
rect 106 62 108 66
rect 116 64 118 69
rect 126 64 128 69
rect 26 40 28 44
rect 36 40 38 51
rect 46 48 48 51
rect 66 48 68 51
rect 46 46 52 48
rect 46 44 48 46
rect 50 44 52 46
rect 46 42 52 44
rect 62 46 68 48
rect 62 44 64 46
rect 66 44 68 46
rect 62 42 68 44
rect 26 38 32 40
rect 26 36 28 38
rect 30 36 32 38
rect 26 34 32 36
rect 36 38 42 40
rect 36 36 38 38
rect 40 36 42 38
rect 36 34 42 36
rect 26 29 28 34
rect 39 29 41 34
rect 46 29 48 42
rect 66 29 68 42
rect 76 40 78 51
rect 86 40 88 44
rect 72 38 78 40
rect 72 36 74 38
rect 76 36 78 38
rect 72 34 78 36
rect 82 38 88 40
rect 82 36 84 38
rect 86 36 88 38
rect 82 34 88 36
rect 73 29 75 34
rect 86 29 88 34
rect 106 40 108 44
rect 116 40 118 51
rect 126 48 128 51
rect 126 46 132 48
rect 126 44 128 46
rect 130 44 132 46
rect 126 42 132 44
rect 140 46 146 48
rect 140 44 142 46
rect 144 44 146 46
rect 191 71 193 75
rect 171 62 173 66
rect 181 62 183 66
rect 140 42 146 44
rect 106 38 112 40
rect 106 36 108 38
rect 110 36 112 38
rect 106 34 112 36
rect 116 38 122 40
rect 116 36 118 38
rect 120 36 122 38
rect 116 34 122 36
rect 106 29 108 34
rect 119 29 121 34
rect 126 29 128 42
rect 144 41 146 42
rect 155 41 157 44
rect 171 41 173 44
rect 144 39 157 41
rect 163 39 173 41
rect 181 40 183 44
rect 191 41 193 44
rect 147 31 149 39
rect 163 35 165 39
rect 156 33 165 35
rect 177 38 183 40
rect 177 36 179 38
rect 181 36 183 38
rect 177 34 183 36
rect 187 39 193 41
rect 187 37 189 39
rect 191 37 193 39
rect 187 35 193 37
rect 156 31 158 33
rect 160 31 165 33
rect 26 16 28 20
rect 39 13 41 18
rect 46 13 48 18
rect 66 13 68 18
rect 73 13 75 18
rect 86 16 88 20
rect 106 16 108 20
rect 156 29 165 31
rect 181 31 183 34
rect 163 26 165 29
rect 173 26 175 30
rect 181 29 185 31
rect 183 26 185 29
rect 190 26 192 35
rect 147 19 149 22
rect 119 13 121 18
rect 126 13 128 18
rect 147 17 152 19
rect 150 9 152 17
rect 163 13 165 17
rect 173 9 175 17
rect 183 9 185 14
rect 190 9 192 14
rect 150 7 175 9
<< ndif >>
rect 37 144 44 146
rect 37 142 40 144
rect 42 142 44 144
rect 37 136 44 142
rect 77 144 84 146
rect 77 142 80 144
rect 82 142 84 144
rect 19 134 26 136
rect 19 132 21 134
rect 23 132 26 134
rect 19 130 26 132
rect 21 125 26 130
rect 28 125 33 136
rect 35 134 44 136
rect 77 136 84 142
rect 106 144 112 146
rect 106 142 108 144
rect 110 142 112 144
rect 106 140 112 142
rect 59 134 66 136
rect 35 125 46 134
rect 48 132 55 134
rect 48 130 51 132
rect 53 130 55 132
rect 59 132 61 134
rect 63 132 66 134
rect 59 130 66 132
rect 48 128 55 130
rect 48 125 53 128
rect 61 125 66 130
rect 68 125 73 136
rect 75 134 84 136
rect 75 125 86 134
rect 88 132 95 134
rect 88 130 91 132
rect 93 130 95 132
rect 88 128 95 130
rect 106 128 114 140
rect 116 128 121 140
rect 123 137 128 140
rect 189 144 196 146
rect 189 142 192 144
rect 194 142 196 144
rect 123 134 131 137
rect 123 132 126 134
rect 128 132 131 134
rect 123 128 131 132
rect 133 132 141 137
rect 133 130 136 132
rect 138 130 141 132
rect 133 128 141 130
rect 143 135 152 137
rect 189 136 196 142
rect 143 133 148 135
rect 150 133 152 135
rect 143 132 152 133
rect 171 134 178 136
rect 171 132 173 134
rect 175 132 178 134
rect 143 128 157 132
rect 88 125 93 128
rect 152 123 157 128
rect 159 129 164 132
rect 171 130 178 132
rect 159 127 166 129
rect 159 125 162 127
rect 164 125 166 127
rect 173 125 178 130
rect 180 125 185 136
rect 187 134 196 136
rect 187 125 198 134
rect 200 132 207 134
rect 200 130 203 132
rect 205 130 207 132
rect 200 128 207 130
rect 200 125 205 128
rect 159 123 166 125
rect 140 29 147 31
rect 21 26 26 29
rect 19 24 26 26
rect 19 22 21 24
rect 23 22 26 24
rect 19 20 26 22
rect 28 20 39 29
rect 30 18 39 20
rect 41 18 46 29
rect 48 24 53 29
rect 61 24 66 29
rect 48 22 55 24
rect 48 20 51 22
rect 53 20 55 22
rect 48 18 55 20
rect 59 22 66 24
rect 59 20 61 22
rect 63 20 66 22
rect 59 18 66 20
rect 68 18 73 29
rect 75 20 86 29
rect 88 26 93 29
rect 101 26 106 29
rect 88 24 95 26
rect 88 22 91 24
rect 93 22 95 24
rect 88 20 95 22
rect 99 24 106 26
rect 99 22 101 24
rect 103 22 106 24
rect 99 20 106 22
rect 108 20 119 29
rect 75 18 84 20
rect 30 12 37 18
rect 30 10 32 12
rect 34 10 37 12
rect 30 8 37 10
rect 77 12 84 18
rect 110 18 119 20
rect 121 18 126 29
rect 128 24 133 29
rect 140 27 142 29
rect 144 27 147 29
rect 140 25 147 27
rect 128 22 135 24
rect 142 22 147 25
rect 149 26 154 31
rect 149 22 163 26
rect 128 20 131 22
rect 133 20 135 22
rect 128 18 135 20
rect 154 21 163 22
rect 154 19 156 21
rect 158 19 163 21
rect 77 10 80 12
rect 82 10 84 12
rect 77 8 84 10
rect 110 12 117 18
rect 154 17 163 19
rect 165 24 173 26
rect 165 22 168 24
rect 170 22 173 24
rect 165 17 173 22
rect 175 22 183 26
rect 175 20 178 22
rect 180 20 183 22
rect 175 17 183 20
rect 110 10 112 12
rect 114 10 117 12
rect 110 8 117 10
rect 178 14 183 17
rect 185 14 190 26
rect 192 14 200 26
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
<< pdif >>
rect 40 103 46 110
rect 19 94 26 103
rect 19 92 21 94
rect 23 92 26 94
rect 19 90 26 92
rect 28 101 36 103
rect 28 99 31 101
rect 33 99 36 101
rect 28 94 36 99
rect 28 92 31 94
rect 33 92 36 94
rect 28 90 36 92
rect 38 96 46 103
rect 38 94 41 96
rect 43 94 46 96
rect 38 92 46 94
rect 48 108 55 110
rect 48 106 51 108
rect 53 106 55 108
rect 48 101 55 106
rect 80 103 86 110
rect 48 99 51 101
rect 53 99 55 101
rect 48 97 55 99
rect 48 92 53 97
rect 59 94 66 103
rect 59 92 61 94
rect 63 92 66 94
rect 38 90 44 92
rect 59 90 66 92
rect 68 101 76 103
rect 68 99 71 101
rect 73 99 76 101
rect 68 94 76 99
rect 68 92 71 94
rect 73 92 76 94
rect 68 90 76 92
rect 78 96 86 103
rect 78 94 81 96
rect 83 94 86 96
rect 78 92 86 94
rect 88 108 95 110
rect 88 106 91 108
rect 93 106 95 108
rect 88 101 95 106
rect 88 99 91 101
rect 93 99 95 101
rect 88 97 95 99
rect 88 92 93 97
rect 108 95 113 110
rect 106 93 113 95
rect 78 90 84 92
rect 106 91 108 93
rect 110 91 113 93
rect 106 89 113 91
rect 108 83 113 89
rect 115 101 123 110
rect 115 99 118 101
rect 120 99 123 101
rect 115 92 123 99
rect 125 108 133 110
rect 125 106 128 108
rect 130 106 133 108
rect 125 101 133 106
rect 125 99 128 101
rect 130 99 133 101
rect 125 92 133 99
rect 135 94 149 110
rect 135 92 144 94
rect 146 92 149 94
rect 115 83 120 92
rect 137 87 149 92
rect 137 85 144 87
rect 146 85 149 87
rect 137 83 149 85
rect 151 108 158 110
rect 151 106 154 108
rect 156 106 158 108
rect 151 104 158 106
rect 151 83 156 104
rect 192 103 198 110
rect 171 94 178 103
rect 171 92 173 94
rect 175 92 178 94
rect 171 90 178 92
rect 180 101 188 103
rect 180 99 183 101
rect 185 99 188 101
rect 180 94 188 99
rect 180 92 183 94
rect 185 92 188 94
rect 180 90 188 92
rect 190 96 198 103
rect 190 94 193 96
rect 195 94 198 96
rect 190 92 198 94
rect 200 108 207 110
rect 200 106 203 108
rect 205 106 207 108
rect 200 101 207 106
rect 200 99 203 101
rect 205 99 207 101
rect 200 97 207 99
rect 200 92 205 97
rect 190 90 196 92
rect 30 62 36 64
rect 21 57 26 62
rect 19 55 26 57
rect 19 53 21 55
rect 23 53 26 55
rect 19 48 26 53
rect 19 46 21 48
rect 23 46 26 48
rect 19 44 26 46
rect 28 60 36 62
rect 28 58 31 60
rect 33 58 36 60
rect 28 51 36 58
rect 38 62 46 64
rect 38 60 41 62
rect 43 60 46 62
rect 38 55 46 60
rect 38 53 41 55
rect 43 53 46 55
rect 38 51 46 53
rect 48 62 55 64
rect 48 60 51 62
rect 53 60 55 62
rect 48 51 55 60
rect 59 62 66 64
rect 59 60 61 62
rect 63 60 66 62
rect 59 51 66 60
rect 68 62 76 64
rect 68 60 71 62
rect 73 60 76 62
rect 68 55 76 60
rect 68 53 71 55
rect 73 53 76 55
rect 68 51 76 53
rect 78 62 84 64
rect 110 62 116 64
rect 78 60 86 62
rect 78 58 81 60
rect 83 58 86 60
rect 78 51 86 58
rect 28 44 34 51
rect 80 44 86 51
rect 88 57 93 62
rect 101 57 106 62
rect 88 55 95 57
rect 88 53 91 55
rect 93 53 95 55
rect 88 48 95 53
rect 88 46 91 48
rect 93 46 95 48
rect 88 44 95 46
rect 99 55 106 57
rect 99 53 101 55
rect 103 53 106 55
rect 99 48 106 53
rect 99 46 101 48
rect 103 46 106 48
rect 99 44 106 46
rect 108 60 116 62
rect 108 58 111 60
rect 113 58 116 60
rect 108 51 116 58
rect 118 62 126 64
rect 118 60 121 62
rect 123 60 126 62
rect 118 55 126 60
rect 118 53 121 55
rect 123 53 126 55
rect 118 51 126 53
rect 128 62 135 64
rect 128 60 131 62
rect 133 60 135 62
rect 128 51 135 60
rect 108 44 114 51
rect 150 50 155 71
rect 148 48 155 50
rect 148 46 150 48
rect 152 46 155 48
rect 148 44 155 46
rect 157 69 169 71
rect 157 67 160 69
rect 162 67 169 69
rect 157 62 169 67
rect 186 62 191 71
rect 157 60 160 62
rect 162 60 171 62
rect 157 44 171 60
rect 173 55 181 62
rect 173 53 176 55
rect 178 53 181 55
rect 173 48 181 53
rect 173 46 176 48
rect 178 46 181 48
rect 173 44 181 46
rect 183 55 191 62
rect 183 53 186 55
rect 188 53 191 55
rect 183 44 191 53
rect 193 65 198 71
rect 193 63 200 65
rect 193 61 196 63
rect 198 61 200 63
rect 193 59 200 61
rect 193 44 198 59
<< alu1 >>
rect 9 144 207 149
rect 9 142 40 144
rect 42 142 50 144
rect 52 142 80 144
rect 82 142 90 144
rect 92 142 108 144
rect 110 142 161 144
rect 163 142 192 144
rect 194 142 202 144
rect 204 142 207 144
rect 9 141 207 142
rect 26 119 31 128
rect 43 132 55 136
rect 43 130 51 132
rect 53 130 55 132
rect 51 127 55 130
rect 26 118 40 119
rect 26 116 34 118
rect 36 116 37 118
rect 39 116 40 118
rect 26 115 40 116
rect 19 110 32 111
rect 19 108 24 110
rect 26 108 32 110
rect 19 107 32 108
rect 19 102 23 107
rect 51 125 52 127
rect 54 125 55 127
rect 51 110 55 125
rect 66 119 71 128
rect 83 132 95 136
rect 83 130 91 132
rect 93 130 95 132
rect 66 118 80 119
rect 66 116 74 118
rect 76 116 77 118
rect 79 116 80 118
rect 66 115 80 116
rect 19 100 20 102
rect 22 100 23 102
rect 19 98 23 100
rect 50 108 55 110
rect 50 106 51 108
rect 53 106 55 108
rect 50 101 55 106
rect 50 99 51 101
rect 53 99 55 101
rect 50 97 55 99
rect 59 110 72 111
rect 59 108 64 110
rect 66 108 72 110
rect 59 107 72 108
rect 59 103 63 107
rect 91 110 95 130
rect 59 101 60 103
rect 62 101 63 103
rect 59 98 63 101
rect 90 108 95 110
rect 90 106 91 108
rect 93 106 95 108
rect 90 104 95 106
rect 90 102 91 104
rect 93 102 95 104
rect 90 101 95 102
rect 90 99 91 101
rect 93 99 95 101
rect 90 97 95 99
rect 106 134 130 135
rect 106 132 126 134
rect 128 132 130 134
rect 106 131 130 132
rect 106 103 110 131
rect 145 127 158 128
rect 145 125 153 127
rect 155 125 158 127
rect 145 123 158 125
rect 145 121 146 123
rect 148 122 158 123
rect 148 121 150 122
rect 106 101 122 103
rect 106 99 118 101
rect 120 99 122 101
rect 106 98 122 99
rect 145 114 150 121
rect 178 127 183 128
rect 178 125 180 127
rect 182 125 183 127
rect 178 119 183 125
rect 195 132 207 136
rect 195 130 203 132
rect 205 130 207 132
rect 178 118 192 119
rect 178 116 186 118
rect 188 116 192 118
rect 178 115 192 116
rect 161 111 166 112
rect 161 110 167 111
rect 171 110 184 111
rect 161 108 162 110
rect 164 108 176 110
rect 178 108 184 110
rect 161 107 184 108
rect 161 105 175 107
rect 161 96 166 105
rect 171 104 175 105
rect 203 115 207 130
rect 203 113 204 115
rect 206 113 207 115
rect 203 110 207 113
rect 171 102 172 104
rect 174 102 175 104
rect 171 98 175 102
rect 202 108 207 110
rect 202 106 203 108
rect 205 106 207 108
rect 202 101 207 106
rect 154 90 166 96
rect 202 99 203 101
rect 205 99 207 101
rect 202 97 207 99
rect 18 84 207 85
rect 18 82 50 84
rect 52 82 90 84
rect 92 82 128 84
rect 130 82 202 84
rect 204 82 207 84
rect 18 72 207 82
rect 18 70 22 72
rect 24 70 90 72
rect 92 70 102 72
rect 104 70 176 72
rect 178 70 207 72
rect 18 69 207 70
rect 19 55 24 57
rect 19 53 21 55
rect 23 53 24 55
rect 19 48 24 53
rect 19 46 21 48
rect 23 46 24 48
rect 19 44 24 46
rect 51 55 55 56
rect 51 53 52 55
rect 54 53 55 55
rect 19 24 23 44
rect 51 47 55 53
rect 42 46 55 47
rect 42 44 48 46
rect 50 44 55 46
rect 42 43 55 44
rect 59 47 63 56
rect 90 55 95 57
rect 59 46 72 47
rect 59 44 60 46
rect 62 44 64 46
rect 66 44 72 46
rect 59 43 72 44
rect 34 38 48 39
rect 34 36 35 38
rect 37 36 38 38
rect 40 36 48 38
rect 34 35 48 36
rect 19 22 21 24
rect 23 22 31 24
rect 19 18 31 22
rect 43 26 48 35
rect 66 38 80 39
rect 66 36 74 38
rect 76 36 77 38
rect 79 36 80 38
rect 66 35 80 36
rect 90 53 91 55
rect 93 53 95 55
rect 90 48 95 53
rect 90 46 91 48
rect 93 46 95 48
rect 90 44 95 46
rect 66 26 71 35
rect 91 29 95 44
rect 91 27 92 29
rect 94 27 95 29
rect 91 24 95 27
rect 83 22 91 24
rect 93 22 95 24
rect 83 18 95 22
rect 99 55 104 57
rect 99 53 101 55
rect 103 53 104 55
rect 140 62 152 64
rect 140 60 148 62
rect 150 60 152 62
rect 140 58 152 60
rect 99 48 104 53
rect 99 46 101 48
rect 103 46 104 48
rect 99 44 104 46
rect 99 24 103 44
rect 131 49 135 56
rect 140 49 145 58
rect 131 47 145 49
rect 122 46 145 47
rect 122 44 128 46
rect 130 44 142 46
rect 144 44 145 46
rect 122 43 135 44
rect 139 43 145 44
rect 140 42 145 43
rect 114 38 128 39
rect 114 36 118 38
rect 120 36 128 38
rect 114 35 128 36
rect 99 22 101 24
rect 103 22 111 24
rect 99 18 111 22
rect 123 29 128 35
rect 123 27 124 29
rect 126 27 128 29
rect 123 26 128 27
rect 156 33 161 40
rect 184 55 200 56
rect 184 53 186 55
rect 188 53 200 55
rect 184 51 200 53
rect 156 32 158 33
rect 148 31 158 32
rect 160 31 161 33
rect 148 29 161 31
rect 148 27 151 29
rect 153 27 161 29
rect 148 26 161 27
rect 196 23 200 51
rect 176 22 200 23
rect 176 20 178 22
rect 180 20 200 22
rect 176 19 200 20
rect 9 12 204 13
rect 9 10 22 12
rect 24 10 32 12
rect 34 10 80 12
rect 82 10 90 12
rect 92 10 102 12
rect 104 10 112 12
rect 114 10 143 12
rect 145 10 196 12
rect 198 10 204 12
rect 9 5 204 10
<< alu2 >>
rect 51 127 183 128
rect 51 125 52 127
rect 54 125 153 127
rect 155 125 180 127
rect 182 125 183 127
rect 51 124 183 125
rect 34 118 40 119
rect 34 116 37 118
rect 39 116 40 118
rect 11 102 23 103
rect 11 100 20 102
rect 22 100 23 102
rect 11 98 23 100
rect 11 25 16 98
rect 34 38 40 116
rect 76 118 80 119
rect 76 116 77 118
rect 79 116 80 118
rect 59 103 63 104
rect 59 101 60 103
rect 62 101 63 103
rect 59 77 63 101
rect 51 73 63 77
rect 51 55 55 73
rect 51 53 52 55
rect 54 53 55 55
rect 51 52 55 53
rect 34 36 35 38
rect 37 36 40 38
rect 34 35 40 36
rect 59 46 63 47
rect 59 44 60 46
rect 62 44 63 46
rect 59 25 63 44
rect 76 38 80 116
rect 203 115 207 119
rect 203 113 204 115
rect 206 113 207 115
rect 90 104 175 105
rect 90 102 91 104
rect 93 102 172 104
rect 174 102 175 104
rect 90 101 175 102
rect 203 78 207 113
rect 147 73 207 78
rect 147 62 152 73
rect 147 60 148 62
rect 150 60 152 62
rect 147 58 152 60
rect 76 36 77 38
rect 79 36 80 38
rect 76 35 80 36
rect 91 29 156 30
rect 91 27 92 29
rect 94 27 124 29
rect 126 27 151 29
rect 153 27 156 29
rect 91 26 156 27
rect 91 25 129 26
rect 11 21 63 25
<< ptie >>
rect 48 144 54 146
rect 48 142 50 144
rect 52 142 54 144
rect 48 140 54 142
rect 88 144 94 146
rect 88 142 90 144
rect 92 142 94 144
rect 88 140 94 142
rect 159 144 165 146
rect 159 142 161 144
rect 163 142 165 144
rect 159 140 165 142
rect 200 144 206 146
rect 200 142 202 144
rect 204 142 206 144
rect 200 140 206 142
rect 20 12 26 14
rect 20 10 22 12
rect 24 10 26 12
rect 20 8 26 10
rect 88 12 94 14
rect 88 10 90 12
rect 92 10 94 12
rect 88 8 94 10
rect 100 12 106 14
rect 100 10 102 12
rect 104 10 106 12
rect 100 8 106 10
rect 141 12 147 14
rect 141 10 143 12
rect 145 10 147 12
rect 141 8 147 10
<< ntie >>
rect 48 84 54 86
rect 48 82 50 84
rect 52 82 54 84
rect 48 80 54 82
rect 88 84 94 86
rect 88 82 90 84
rect 92 82 94 84
rect 126 84 132 86
rect 88 80 94 82
rect 126 82 128 84
rect 130 82 132 84
rect 200 84 206 86
rect 126 80 132 82
rect 200 82 202 84
rect 204 82 206 84
rect 200 80 206 82
rect 20 72 26 74
rect 20 70 22 72
rect 24 70 26 72
rect 20 68 26 70
rect 88 72 94 74
rect 88 70 90 72
rect 92 70 94 72
rect 88 68 94 70
rect 100 72 106 74
rect 100 70 102 72
rect 104 70 106 72
rect 174 72 180 74
rect 100 68 106 70
rect 174 70 176 72
rect 178 70 180 72
rect 174 68 180 70
<< nmos >>
rect 26 125 28 136
rect 33 125 35 136
rect 46 125 48 134
rect 66 125 68 136
rect 73 125 75 136
rect 86 125 88 134
rect 114 128 116 140
rect 121 128 123 140
rect 131 128 133 137
rect 141 128 143 137
rect 157 123 159 132
rect 178 125 180 136
rect 185 125 187 136
rect 198 125 200 134
rect 26 20 28 29
rect 39 18 41 29
rect 46 18 48 29
rect 66 18 68 29
rect 73 18 75 29
rect 86 20 88 29
rect 106 20 108 29
rect 119 18 121 29
rect 126 18 128 29
rect 147 22 149 31
rect 163 17 165 26
rect 173 17 175 26
rect 183 14 185 26
rect 190 14 192 26
<< pmos >>
rect 26 90 28 103
rect 36 90 38 103
rect 46 92 48 110
rect 66 90 68 103
rect 76 90 78 103
rect 86 92 88 110
rect 113 83 115 110
rect 123 92 125 110
rect 133 92 135 110
rect 149 83 151 110
rect 178 90 180 103
rect 188 90 190 103
rect 198 92 200 110
rect 26 44 28 62
rect 36 51 38 64
rect 46 51 48 64
rect 66 51 68 64
rect 76 51 78 64
rect 86 44 88 62
rect 106 44 108 62
rect 116 51 118 64
rect 126 51 128 64
rect 155 44 157 71
rect 171 44 173 62
rect 181 44 183 62
rect 191 44 193 71
<< polyct0 >>
rect 44 116 46 118
rect 84 116 86 118
rect 115 115 117 117
rect 125 116 127 118
rect 196 116 198 118
rect 28 36 30 38
rect 84 36 86 38
rect 108 36 110 38
rect 179 36 181 38
rect 189 37 191 39
<< polyct1 >>
rect 34 116 36 118
rect 24 108 26 110
rect 74 116 76 118
rect 146 121 148 123
rect 64 108 66 110
rect 186 116 188 118
rect 162 108 164 110
rect 176 108 178 110
rect 48 44 50 46
rect 64 44 66 46
rect 38 36 40 38
rect 74 36 76 38
rect 128 44 130 46
rect 142 44 144 46
rect 118 36 120 38
rect 158 31 160 33
<< ndifct0 >>
rect 21 132 23 134
rect 61 132 63 134
rect 136 130 138 132
rect 148 133 150 135
rect 173 132 175 134
rect 162 125 164 127
rect 51 20 53 22
rect 61 20 63 22
rect 142 27 144 29
rect 131 20 133 22
rect 156 19 158 21
rect 168 22 170 24
<< ndifct1 >>
rect 40 142 42 144
rect 80 142 82 144
rect 108 142 110 144
rect 51 130 53 132
rect 91 130 93 132
rect 192 142 194 144
rect 126 132 128 134
rect 203 130 205 132
rect 21 22 23 24
rect 91 22 93 24
rect 101 22 103 24
rect 32 10 34 12
rect 80 10 82 12
rect 178 20 180 22
rect 112 10 114 12
rect 196 10 198 12
<< ntiect1 >>
rect 50 82 52 84
rect 90 82 92 84
rect 128 82 130 84
rect 202 82 204 84
rect 22 70 24 72
rect 90 70 92 72
rect 102 70 104 72
rect 176 70 178 72
<< ptiect1 >>
rect 50 142 52 144
rect 90 142 92 144
rect 161 142 163 144
rect 202 142 204 144
rect 22 10 24 12
rect 90 10 92 12
rect 102 10 104 12
rect 143 10 145 12
<< pdifct0 >>
rect 21 92 23 94
rect 31 99 33 101
rect 31 92 33 94
rect 41 94 43 96
rect 61 92 63 94
rect 71 99 73 101
rect 71 92 73 94
rect 81 94 83 96
rect 108 91 110 93
rect 128 106 130 108
rect 128 99 130 101
rect 144 92 146 94
rect 144 85 146 87
rect 154 106 156 108
rect 173 92 175 94
rect 183 99 185 101
rect 183 92 185 94
rect 193 94 195 96
rect 31 58 33 60
rect 41 60 43 62
rect 41 53 43 55
rect 51 60 53 62
rect 61 60 63 62
rect 71 60 73 62
rect 71 53 73 55
rect 81 58 83 60
rect 111 58 113 60
rect 121 60 123 62
rect 121 53 123 55
rect 131 60 133 62
rect 150 46 152 48
rect 160 67 162 69
rect 160 60 162 62
rect 176 53 178 55
rect 176 46 178 48
rect 196 61 198 63
<< pdifct1 >>
rect 51 106 53 108
rect 51 99 53 101
rect 91 106 93 108
rect 91 99 93 101
rect 118 99 120 101
rect 203 106 205 108
rect 203 99 205 101
rect 21 53 23 55
rect 21 46 23 48
rect 91 53 93 55
rect 91 46 93 48
rect 101 53 103 55
rect 101 46 103 48
rect 186 53 188 55
<< alu0 >>
rect 19 134 39 135
rect 19 132 21 134
rect 23 132 39 134
rect 19 131 39 132
rect 35 127 39 131
rect 59 134 79 135
rect 59 132 61 134
rect 63 132 79 134
rect 59 131 79 132
rect 50 128 51 130
rect 35 123 47 127
rect 43 118 47 123
rect 43 116 44 118
rect 46 116 47 118
rect 43 104 47 116
rect 75 127 79 131
rect 146 135 152 141
rect 90 128 91 130
rect 75 123 87 127
rect 83 118 87 123
rect 83 116 84 118
rect 86 116 87 118
rect 30 101 47 104
rect 30 99 31 101
rect 33 100 47 101
rect 33 99 34 100
rect 19 94 25 95
rect 19 92 21 94
rect 23 92 25 94
rect 19 85 25 92
rect 30 94 34 99
rect 83 104 87 116
rect 70 101 87 104
rect 70 99 71 101
rect 73 100 87 101
rect 73 99 74 100
rect 30 92 31 94
rect 33 92 34 94
rect 30 90 34 92
rect 39 96 45 97
rect 39 94 41 96
rect 43 94 45 96
rect 39 85 45 94
rect 59 94 65 95
rect 59 92 61 94
rect 63 92 65 94
rect 59 85 65 92
rect 70 94 74 99
rect 135 132 139 134
rect 146 133 148 135
rect 150 133 152 135
rect 146 132 152 133
rect 171 134 191 135
rect 171 132 173 134
rect 175 132 191 134
rect 135 130 136 132
rect 138 130 139 132
rect 171 131 191 132
rect 135 127 139 130
rect 115 123 139 127
rect 115 119 119 123
rect 161 127 165 129
rect 161 125 162 127
rect 164 125 165 127
rect 114 117 119 119
rect 114 115 115 117
rect 117 115 119 117
rect 123 118 139 119
rect 123 116 125 118
rect 127 116 139 118
rect 123 115 139 116
rect 114 113 119 115
rect 115 111 119 113
rect 115 108 131 111
rect 115 107 128 108
rect 127 106 128 107
rect 130 106 131 108
rect 127 101 131 106
rect 127 99 128 101
rect 130 99 131 101
rect 127 97 131 99
rect 135 109 139 115
rect 161 119 165 125
rect 154 115 165 119
rect 187 127 191 131
rect 202 128 203 130
rect 187 123 199 127
rect 195 118 199 123
rect 195 116 196 118
rect 198 116 199 118
rect 154 109 158 115
rect 135 108 158 109
rect 135 106 154 108
rect 156 106 158 108
rect 135 105 158 106
rect 70 92 71 94
rect 73 92 74 94
rect 70 90 74 92
rect 79 96 85 97
rect 79 94 81 96
rect 83 94 85 96
rect 135 94 139 105
rect 195 104 199 116
rect 182 101 199 104
rect 182 99 183 101
rect 185 100 199 101
rect 185 99 186 100
rect 79 85 85 94
rect 106 93 139 94
rect 106 91 108 93
rect 110 91 139 93
rect 106 90 139 91
rect 143 94 147 96
rect 143 92 144 94
rect 146 92 147 94
rect 143 87 147 92
rect 171 94 177 95
rect 171 92 173 94
rect 175 92 177 94
rect 143 85 144 87
rect 146 85 147 87
rect 171 85 177 92
rect 182 94 186 99
rect 182 92 183 94
rect 185 92 186 94
rect 182 90 186 92
rect 191 96 197 97
rect 191 94 193 96
rect 195 94 197 96
rect 191 85 197 94
rect 29 60 35 69
rect 29 58 31 60
rect 33 58 35 60
rect 29 57 35 58
rect 40 62 44 64
rect 40 60 41 62
rect 43 60 44 62
rect 40 55 44 60
rect 49 62 55 69
rect 49 60 51 62
rect 53 60 55 62
rect 49 59 55 60
rect 59 62 65 69
rect 59 60 61 62
rect 63 60 65 62
rect 59 59 65 60
rect 70 62 74 64
rect 70 60 71 62
rect 73 60 74 62
rect 40 54 41 55
rect 27 53 41 54
rect 43 53 44 55
rect 27 50 44 53
rect 27 38 31 50
rect 70 55 74 60
rect 79 60 85 69
rect 79 58 81 60
rect 83 58 85 60
rect 79 57 85 58
rect 109 60 115 69
rect 109 58 111 60
rect 113 58 115 60
rect 109 57 115 58
rect 120 62 124 64
rect 120 60 121 62
rect 123 60 124 62
rect 70 53 71 55
rect 73 54 74 55
rect 73 53 87 54
rect 70 50 87 53
rect 27 36 28 38
rect 30 36 31 38
rect 27 31 31 36
rect 27 27 39 31
rect 23 24 24 26
rect 35 23 39 27
rect 83 38 87 50
rect 83 36 84 38
rect 86 36 87 38
rect 83 31 87 36
rect 75 27 87 31
rect 75 23 79 27
rect 90 24 91 26
rect 35 22 55 23
rect 35 20 51 22
rect 53 20 55 22
rect 35 19 55 20
rect 59 22 79 23
rect 59 20 61 22
rect 63 20 79 22
rect 59 19 79 20
rect 120 55 124 60
rect 129 62 135 69
rect 159 67 160 69
rect 162 67 163 69
rect 129 60 131 62
rect 133 60 135 62
rect 129 59 135 60
rect 159 62 163 67
rect 159 60 160 62
rect 162 60 163 62
rect 159 58 163 60
rect 167 63 200 64
rect 167 61 196 63
rect 198 61 200 63
rect 167 60 200 61
rect 120 54 121 55
rect 107 53 121 54
rect 123 53 124 55
rect 107 50 124 53
rect 107 38 111 50
rect 167 49 171 60
rect 148 48 171 49
rect 148 46 150 48
rect 152 46 171 48
rect 148 45 171 46
rect 148 39 152 45
rect 107 36 108 38
rect 110 36 111 38
rect 107 31 111 36
rect 107 27 119 31
rect 103 24 104 26
rect 115 23 119 27
rect 141 35 152 39
rect 141 29 145 35
rect 167 39 171 45
rect 175 55 179 57
rect 175 53 176 55
rect 178 53 179 55
rect 175 48 179 53
rect 175 46 176 48
rect 178 47 179 48
rect 178 46 191 47
rect 175 43 191 46
rect 187 41 191 43
rect 187 39 192 41
rect 167 38 183 39
rect 167 36 179 38
rect 181 36 183 38
rect 167 35 183 36
rect 187 37 189 39
rect 191 37 192 39
rect 187 35 192 37
rect 141 27 142 29
rect 144 27 145 29
rect 141 25 145 27
rect 187 31 191 35
rect 167 27 191 31
rect 167 24 171 27
rect 115 22 135 23
rect 167 22 168 24
rect 170 22 171 24
rect 115 20 131 22
rect 133 20 135 22
rect 115 19 135 20
rect 154 21 160 22
rect 154 19 156 21
rect 158 19 160 21
rect 167 20 171 22
rect 154 13 160 19
<< via1 >>
rect 37 116 39 118
rect 52 125 54 127
rect 77 116 79 118
rect 20 100 22 102
rect 60 101 62 103
rect 91 102 93 104
rect 153 125 155 127
rect 180 125 182 127
rect 204 113 206 115
rect 172 102 174 104
rect 52 53 54 55
rect 60 44 62 46
rect 35 36 37 38
rect 77 36 79 38
rect 92 27 94 29
rect 148 60 150 62
rect 124 27 126 29
rect 151 27 153 29
<< labels >>
rlabel alu1 141 73 141 73 1 Vdd
rlabel alu1 117 73 117 73 6 vdd
rlabel alu1 139 8 139 8 1 Vss
rlabel alu1 37 9 37 9 6 vss
rlabel alu1 37 73 37 73 6 vdd
rlabel alu1 45 31 45 31 1 a0
rlabel alu1 53 53 53 53 1 b0
rlabel alu1 61 53 61 53 1 b1
rlabel alu1 69 32 69 32 1 a1
rlabel alu1 77 9 77 9 4 vss
rlabel alu1 77 73 77 73 4 vdd
rlabel alu1 167 146 167 146 5 Vss
rlabel alu1 189 81 189 81 2 vdd
rlabel alu1 165 81 165 81 5 Vdd
rlabel alu1 37 81 37 81 2 vdd
rlabel alu1 37 145 37 145 2 vss
rlabel alu1 77 145 77 145 2 vss
rlabel alu1 77 81 77 81 2 vdd
rlabel alu1 69 109 69 109 1 b0
rlabel alu1 69 121 69 121 1 a1
rlabel alu1 29 123 29 123 1 a0
rlabel via1 21 101 21 101 1 b1
rlabel alu1 21 37 21 37 1 r0
rlabel alu1 108 114 108 114 1 r1
rlabel alu1 198 40 198 40 1 p02
rlabel alu1 101 35 101 35 1 p03
<< end >>
