magic
tech scmos
timestamp 1608969680
<< ab >>
rect 191 340 239 348
rect 200 275 239 340
rect 241 275 277 348
rect 200 212 237 275
rect 191 204 237 212
rect 239 204 277 275
rect 279 340 284 348
rect 279 284 281 340
rect 279 275 284 284
rect 286 275 349 348
rect 351 340 455 348
rect 351 316 389 340
rect 351 275 398 316
rect 279 204 319 275
rect 321 204 384 275
rect 389 236 398 275
rect 416 275 455 340
rect 457 275 493 348
rect 416 212 453 275
rect 385 204 453 212
rect 455 204 493 275
rect 495 340 500 348
rect 495 284 497 340
rect 495 275 500 284
rect 502 275 565 348
rect 567 340 660 348
rect 567 316 605 340
rect 567 284 614 316
rect 621 284 660 340
rect 567 275 660 284
rect 662 275 698 348
rect 495 204 535 275
rect 537 204 600 275
rect 605 268 658 275
rect 605 236 614 268
rect 621 212 658 268
rect 602 204 658 212
rect 660 204 698 275
rect 700 340 705 348
rect 700 284 702 340
rect 700 275 705 284
rect 707 275 770 348
rect 772 340 879 348
rect 772 316 810 340
rect 772 275 819 316
rect 700 204 740 275
rect 742 204 805 275
rect 810 236 819 275
rect 840 275 879 340
rect 881 275 917 348
rect 840 212 877 275
rect 807 204 877 212
rect 879 204 917 275
rect 919 340 924 348
rect 919 284 921 340
rect 919 275 924 284
rect 926 275 989 348
rect 991 316 1029 348
rect 991 275 1038 316
rect 919 204 959 275
rect 961 204 1024 275
rect 1029 236 1038 275
rect 1043 204 1083 276
rect 1085 204 1148 276
rect 149 132 229 204
rect 231 132 334 204
rect 336 132 479 204
rect 481 132 584 204
rect 586 132 729 204
rect 731 132 834 204
rect 836 132 979 204
rect 981 132 1084 204
rect 1086 132 1149 204
rect 148 60 228 132
rect 230 60 333 132
rect 335 60 478 132
rect 480 60 583 132
rect 585 60 728 132
rect 730 60 833 132
rect 835 60 978 132
rect 980 89 1083 132
rect 1085 89 1148 132
rect 980 87 1148 89
rect 980 60 1083 87
rect 1085 60 1148 87
rect 147 -12 227 60
rect 229 52 332 60
rect 229 43 242 52
rect 244 43 332 52
rect 229 -12 332 43
rect 334 -12 477 60
rect 479 -12 582 60
rect 584 -12 727 60
rect 729 -12 832 60
rect 834 -12 977 60
rect 979 33 1082 60
rect 1084 33 1147 60
rect 979 31 1147 33
rect 979 -12 1082 31
rect 1084 -12 1147 31
<< nwell >>
rect 182 281 1038 316
rect 182 236 1153 281
rect 144 137 1154 172
rect 143 127 1154 137
rect 143 92 1153 127
rect 142 -17 1152 28
<< pwell >>
rect 182 316 1038 353
rect 182 209 1153 236
rect 144 172 1154 209
rect 143 65 1153 92
rect 142 55 1153 65
rect 142 28 1152 55
<< poly >>
rect 208 335 210 340
rect 215 335 217 340
rect 228 333 230 337
rect 248 335 250 340
rect 255 335 257 340
rect 313 344 338 346
rect 296 339 298 344
rect 303 339 305 344
rect 268 333 270 337
rect 313 336 315 344
rect 323 336 325 340
rect 336 336 338 344
rect 336 334 341 336
rect 360 335 362 340
rect 367 335 369 340
rect 339 331 341 334
rect 208 311 210 324
rect 215 319 217 324
rect 228 319 230 324
rect 214 317 220 319
rect 214 315 216 317
rect 218 315 220 317
rect 214 313 220 315
rect 224 317 230 319
rect 224 315 226 317
rect 228 315 230 317
rect 224 313 230 315
rect 204 309 210 311
rect 204 307 206 309
rect 208 307 210 309
rect 204 305 210 307
rect 208 302 210 305
rect 218 302 220 313
rect 228 309 230 313
rect 248 311 250 324
rect 255 319 257 324
rect 268 319 270 324
rect 254 317 260 319
rect 254 315 256 317
rect 258 315 260 317
rect 254 313 260 315
rect 264 317 270 319
rect 296 318 298 327
rect 303 324 305 327
rect 303 322 307 324
rect 313 323 315 327
rect 323 324 325 327
rect 305 319 307 322
rect 323 322 332 324
rect 380 333 382 337
rect 424 335 426 340
rect 431 335 433 340
rect 444 333 446 337
rect 464 335 466 340
rect 471 335 473 340
rect 529 344 554 346
rect 512 339 514 344
rect 519 339 521 344
rect 484 333 486 337
rect 529 336 531 344
rect 539 336 541 340
rect 552 336 554 344
rect 552 334 557 336
rect 576 335 578 340
rect 583 335 585 340
rect 555 331 557 334
rect 323 320 328 322
rect 330 320 332 322
rect 264 315 266 317
rect 268 315 270 317
rect 264 313 270 315
rect 244 309 250 311
rect 244 307 246 309
rect 248 307 250 309
rect 244 305 250 307
rect 248 302 250 305
rect 258 302 260 313
rect 268 309 270 313
rect 295 316 301 318
rect 295 314 297 316
rect 299 314 301 316
rect 295 312 301 314
rect 305 317 311 319
rect 305 315 307 317
rect 309 315 311 317
rect 305 313 311 315
rect 323 318 332 320
rect 323 314 325 318
rect 339 314 341 322
rect 295 309 297 312
rect 305 309 307 313
rect 315 312 325 314
rect 331 312 344 314
rect 315 309 317 312
rect 331 309 333 312
rect 342 311 344 312
rect 360 311 362 324
rect 367 319 369 324
rect 380 319 382 324
rect 366 317 372 319
rect 366 315 368 317
rect 370 315 372 317
rect 366 313 372 315
rect 376 317 382 319
rect 376 315 378 317
rect 380 315 382 317
rect 376 313 382 315
rect 342 309 348 311
rect 208 284 210 289
rect 218 284 220 289
rect 228 287 230 291
rect 248 284 250 289
rect 258 284 260 289
rect 268 287 270 291
rect 305 287 307 291
rect 315 287 317 291
rect 295 278 297 282
rect 342 307 344 309
rect 346 307 348 309
rect 342 305 348 307
rect 356 309 362 311
rect 356 307 358 309
rect 360 307 362 309
rect 356 305 362 307
rect 360 302 362 305
rect 370 302 372 313
rect 380 309 382 313
rect 424 311 426 324
rect 431 319 433 324
rect 444 319 446 324
rect 430 317 436 319
rect 430 315 432 317
rect 434 315 436 317
rect 430 313 436 315
rect 440 317 446 319
rect 440 315 442 317
rect 444 315 446 317
rect 440 313 446 315
rect 420 309 426 311
rect 420 307 422 309
rect 424 307 426 309
rect 420 305 426 307
rect 424 302 426 305
rect 434 302 436 313
rect 444 309 446 313
rect 464 311 466 324
rect 471 319 473 324
rect 484 319 486 324
rect 470 317 476 319
rect 470 315 472 317
rect 474 315 476 317
rect 470 313 476 315
rect 480 317 486 319
rect 512 318 514 327
rect 519 324 521 327
rect 519 322 523 324
rect 529 323 531 327
rect 539 324 541 327
rect 521 319 523 322
rect 539 322 548 324
rect 596 333 598 337
rect 629 335 631 340
rect 636 335 638 340
rect 649 333 651 337
rect 669 335 671 340
rect 676 335 678 340
rect 734 344 759 346
rect 717 339 719 344
rect 724 339 726 344
rect 689 333 691 337
rect 734 336 736 344
rect 744 336 746 340
rect 757 336 759 344
rect 757 334 762 336
rect 781 335 783 340
rect 788 335 790 340
rect 760 331 762 334
rect 539 320 544 322
rect 546 320 548 322
rect 480 315 482 317
rect 484 315 486 317
rect 480 313 486 315
rect 460 309 466 311
rect 360 284 362 289
rect 370 284 372 289
rect 380 287 382 291
rect 460 307 462 309
rect 464 307 466 309
rect 460 305 466 307
rect 464 302 466 305
rect 474 302 476 313
rect 484 309 486 313
rect 511 316 517 318
rect 511 314 513 316
rect 515 314 517 316
rect 511 312 517 314
rect 521 317 527 319
rect 521 315 523 317
rect 525 315 527 317
rect 521 313 527 315
rect 539 318 548 320
rect 539 314 541 318
rect 555 314 557 322
rect 511 309 513 312
rect 521 309 523 313
rect 531 312 541 314
rect 547 312 560 314
rect 531 309 533 312
rect 547 309 549 312
rect 558 311 560 312
rect 576 311 578 324
rect 583 319 585 324
rect 596 319 598 324
rect 582 317 588 319
rect 582 315 584 317
rect 586 315 588 317
rect 582 313 588 315
rect 592 317 598 319
rect 592 315 594 317
rect 596 315 598 317
rect 592 313 598 315
rect 558 309 564 311
rect 424 284 426 289
rect 434 284 436 289
rect 444 287 446 291
rect 331 278 333 282
rect 464 284 466 289
rect 474 284 476 289
rect 484 287 486 291
rect 521 287 523 291
rect 531 287 533 291
rect 511 278 513 282
rect 558 307 560 309
rect 562 307 564 309
rect 558 305 564 307
rect 572 309 578 311
rect 572 307 574 309
rect 576 307 578 309
rect 572 305 578 307
rect 576 302 578 305
rect 586 302 588 313
rect 596 309 598 313
rect 629 311 631 324
rect 636 319 638 324
rect 649 319 651 324
rect 635 317 641 319
rect 635 315 637 317
rect 639 315 641 317
rect 635 313 641 315
rect 645 317 651 319
rect 645 315 647 317
rect 649 315 651 317
rect 645 313 651 315
rect 625 309 631 311
rect 625 307 627 309
rect 629 307 631 309
rect 625 305 631 307
rect 629 302 631 305
rect 639 302 641 313
rect 649 309 651 313
rect 669 311 671 324
rect 676 319 678 324
rect 689 319 691 324
rect 675 317 681 319
rect 675 315 677 317
rect 679 315 681 317
rect 675 313 681 315
rect 685 317 691 319
rect 717 318 719 327
rect 724 324 726 327
rect 724 322 728 324
rect 734 323 736 327
rect 744 324 746 327
rect 726 319 728 322
rect 744 322 753 324
rect 801 333 803 337
rect 848 335 850 340
rect 855 335 857 340
rect 868 333 870 337
rect 888 335 890 340
rect 895 335 897 340
rect 953 344 978 346
rect 936 339 938 344
rect 943 339 945 344
rect 908 333 910 337
rect 953 336 955 344
rect 963 336 965 340
rect 976 336 978 344
rect 976 334 981 336
rect 1000 335 1002 340
rect 1007 335 1009 340
rect 979 331 981 334
rect 744 320 749 322
rect 751 320 753 322
rect 685 315 687 317
rect 689 315 691 317
rect 685 313 691 315
rect 665 309 671 311
rect 576 284 578 289
rect 586 284 588 289
rect 596 287 598 291
rect 665 307 667 309
rect 669 307 671 309
rect 665 305 671 307
rect 669 302 671 305
rect 679 302 681 313
rect 689 309 691 313
rect 716 316 722 318
rect 716 314 718 316
rect 720 314 722 316
rect 716 312 722 314
rect 726 317 732 319
rect 726 315 728 317
rect 730 315 732 317
rect 726 313 732 315
rect 744 318 753 320
rect 744 314 746 318
rect 760 314 762 322
rect 716 309 718 312
rect 726 309 728 313
rect 736 312 746 314
rect 752 312 765 314
rect 736 309 738 312
rect 752 309 754 312
rect 763 311 765 312
rect 781 311 783 324
rect 788 319 790 324
rect 801 319 803 324
rect 787 317 793 319
rect 787 315 789 317
rect 791 315 793 317
rect 787 313 793 315
rect 797 317 803 319
rect 797 315 799 317
rect 801 315 803 317
rect 797 313 803 315
rect 763 309 769 311
rect 629 284 631 289
rect 639 284 641 289
rect 649 287 651 291
rect 547 278 549 282
rect 669 284 671 289
rect 679 284 681 289
rect 689 287 691 291
rect 726 287 728 291
rect 736 287 738 291
rect 716 278 718 282
rect 763 307 765 309
rect 767 307 769 309
rect 763 305 769 307
rect 777 309 783 311
rect 777 307 779 309
rect 781 307 783 309
rect 777 305 783 307
rect 781 302 783 305
rect 791 302 793 313
rect 801 309 803 313
rect 848 311 850 324
rect 855 319 857 324
rect 868 319 870 324
rect 854 317 860 319
rect 854 315 856 317
rect 858 315 860 317
rect 854 313 860 315
rect 864 317 870 319
rect 864 315 866 317
rect 868 315 870 317
rect 864 313 870 315
rect 844 309 850 311
rect 844 307 846 309
rect 848 307 850 309
rect 844 305 850 307
rect 848 302 850 305
rect 858 302 860 313
rect 868 309 870 313
rect 888 311 890 324
rect 895 319 897 324
rect 908 319 910 324
rect 894 317 900 319
rect 894 315 896 317
rect 898 315 900 317
rect 894 313 900 315
rect 904 317 910 319
rect 936 318 938 327
rect 943 324 945 327
rect 943 322 947 324
rect 953 323 955 327
rect 963 324 965 327
rect 945 319 947 322
rect 963 322 972 324
rect 1020 333 1022 337
rect 963 320 968 322
rect 970 320 972 322
rect 904 315 906 317
rect 908 315 910 317
rect 904 313 910 315
rect 884 309 890 311
rect 781 284 783 289
rect 791 284 793 289
rect 801 287 803 291
rect 884 307 886 309
rect 888 307 890 309
rect 884 305 890 307
rect 888 302 890 305
rect 898 302 900 313
rect 908 309 910 313
rect 935 316 941 318
rect 935 314 937 316
rect 939 314 941 316
rect 935 312 941 314
rect 945 317 951 319
rect 945 315 947 317
rect 949 315 951 317
rect 945 313 951 315
rect 963 318 972 320
rect 963 314 965 318
rect 979 314 981 322
rect 935 309 937 312
rect 945 309 947 313
rect 955 312 965 314
rect 971 312 984 314
rect 955 309 957 312
rect 971 309 973 312
rect 982 311 984 312
rect 1000 311 1002 324
rect 1007 319 1009 324
rect 1020 319 1022 324
rect 1006 317 1012 319
rect 1006 315 1008 317
rect 1010 315 1012 317
rect 1006 313 1012 315
rect 1016 317 1022 319
rect 1016 315 1018 317
rect 1020 315 1022 317
rect 1016 313 1022 315
rect 982 309 988 311
rect 848 284 850 289
rect 858 284 860 289
rect 868 287 870 291
rect 752 278 754 282
rect 888 284 890 289
rect 898 284 900 289
rect 908 287 910 291
rect 945 287 947 291
rect 955 287 957 291
rect 935 278 937 282
rect 982 307 984 309
rect 986 307 988 309
rect 982 305 988 307
rect 996 309 1002 311
rect 996 307 998 309
rect 1000 307 1002 309
rect 996 305 1002 307
rect 1000 302 1002 305
rect 1010 302 1012 313
rect 1020 309 1022 313
rect 1000 284 1002 289
rect 1010 284 1012 289
rect 1020 287 1022 291
rect 971 278 973 282
rect 208 261 210 265
rect 218 263 220 268
rect 228 263 230 268
rect 248 263 250 268
rect 258 263 260 268
rect 337 270 339 274
rect 268 261 270 265
rect 288 261 290 265
rect 298 263 300 268
rect 308 263 310 268
rect 208 239 210 243
rect 218 239 220 250
rect 228 247 230 250
rect 248 247 250 250
rect 228 245 234 247
rect 228 243 230 245
rect 232 243 234 245
rect 228 241 234 243
rect 244 245 250 247
rect 244 243 246 245
rect 248 243 250 245
rect 244 241 250 243
rect 208 237 214 239
rect 208 235 210 237
rect 212 235 214 237
rect 208 233 214 235
rect 218 237 224 239
rect 218 235 220 237
rect 222 235 224 237
rect 218 233 224 235
rect 208 228 210 233
rect 221 228 223 233
rect 228 228 230 241
rect 248 228 250 241
rect 258 239 260 250
rect 268 239 270 243
rect 254 237 260 239
rect 254 235 256 237
rect 258 235 260 237
rect 254 233 260 235
rect 264 237 270 239
rect 264 235 266 237
rect 268 235 270 237
rect 264 233 270 235
rect 255 228 257 233
rect 268 228 270 233
rect 288 239 290 243
rect 298 239 300 250
rect 308 247 310 250
rect 308 245 314 247
rect 308 243 310 245
rect 312 243 314 245
rect 308 241 314 243
rect 322 245 328 247
rect 322 243 324 245
rect 326 243 328 245
rect 373 270 375 274
rect 353 261 355 265
rect 363 261 365 265
rect 424 261 426 265
rect 434 263 436 268
rect 444 263 446 268
rect 464 263 466 268
rect 474 263 476 268
rect 553 270 555 274
rect 484 261 486 265
rect 504 261 506 265
rect 514 263 516 268
rect 524 263 526 268
rect 322 241 328 243
rect 288 237 294 239
rect 288 235 290 237
rect 292 235 294 237
rect 288 233 294 235
rect 298 237 304 239
rect 298 235 300 237
rect 302 235 304 237
rect 298 233 304 235
rect 288 228 290 233
rect 301 228 303 233
rect 308 228 310 241
rect 326 240 328 241
rect 337 240 339 243
rect 353 240 355 243
rect 326 238 339 240
rect 345 238 355 240
rect 363 239 365 243
rect 373 240 375 243
rect 329 230 331 238
rect 345 234 347 238
rect 338 232 347 234
rect 359 237 365 239
rect 359 235 361 237
rect 363 235 365 237
rect 359 233 365 235
rect 369 238 375 240
rect 369 236 371 238
rect 373 236 375 238
rect 369 234 375 236
rect 424 239 426 243
rect 434 239 436 250
rect 444 247 446 250
rect 464 247 466 250
rect 444 245 450 247
rect 444 243 446 245
rect 448 243 450 245
rect 444 241 450 243
rect 460 245 466 247
rect 460 243 462 245
rect 464 243 466 245
rect 460 241 466 243
rect 424 237 430 239
rect 424 235 426 237
rect 428 235 430 237
rect 338 230 340 232
rect 342 230 347 232
rect 208 215 210 219
rect 221 212 223 217
rect 228 212 230 217
rect 248 212 250 217
rect 255 212 257 217
rect 268 215 270 219
rect 288 215 290 219
rect 338 228 347 230
rect 363 230 365 233
rect 345 225 347 228
rect 355 225 357 229
rect 363 228 367 230
rect 365 225 367 228
rect 372 225 374 234
rect 424 233 430 235
rect 434 237 440 239
rect 434 235 436 237
rect 438 235 440 237
rect 434 233 440 235
rect 424 228 426 233
rect 437 228 439 233
rect 444 228 446 241
rect 464 228 466 241
rect 474 239 476 250
rect 484 239 486 243
rect 470 237 476 239
rect 470 235 472 237
rect 474 235 476 237
rect 470 233 476 235
rect 480 237 486 239
rect 480 235 482 237
rect 484 235 486 237
rect 480 233 486 235
rect 471 228 473 233
rect 484 228 486 233
rect 504 239 506 243
rect 514 239 516 250
rect 524 247 526 250
rect 524 245 530 247
rect 524 243 526 245
rect 528 243 530 245
rect 524 241 530 243
rect 538 245 544 247
rect 538 243 540 245
rect 542 243 544 245
rect 589 270 591 274
rect 569 261 571 265
rect 579 261 581 265
rect 629 261 631 265
rect 639 263 641 268
rect 649 263 651 268
rect 669 263 671 268
rect 679 263 681 268
rect 758 270 760 274
rect 689 261 691 265
rect 709 261 711 265
rect 719 263 721 268
rect 729 263 731 268
rect 538 241 544 243
rect 504 237 510 239
rect 504 235 506 237
rect 508 235 510 237
rect 504 233 510 235
rect 514 237 520 239
rect 514 235 516 237
rect 518 235 520 237
rect 514 233 520 235
rect 504 228 506 233
rect 517 228 519 233
rect 524 228 526 241
rect 542 240 544 241
rect 553 240 555 243
rect 569 240 571 243
rect 542 238 555 240
rect 561 238 571 240
rect 579 239 581 243
rect 589 240 591 243
rect 545 230 547 238
rect 561 234 563 238
rect 554 232 563 234
rect 575 237 581 239
rect 575 235 577 237
rect 579 235 581 237
rect 575 233 581 235
rect 585 238 591 240
rect 585 236 587 238
rect 589 236 591 238
rect 585 234 591 236
rect 629 239 631 243
rect 639 239 641 250
rect 649 247 651 250
rect 669 247 671 250
rect 649 245 655 247
rect 649 243 651 245
rect 653 243 655 245
rect 649 241 655 243
rect 665 245 671 247
rect 665 243 667 245
rect 669 243 671 245
rect 665 241 671 243
rect 629 237 635 239
rect 629 235 631 237
rect 633 235 635 237
rect 554 230 556 232
rect 558 230 563 232
rect 329 218 331 221
rect 301 212 303 217
rect 308 212 310 217
rect 329 216 334 218
rect 332 208 334 216
rect 345 212 347 216
rect 355 208 357 216
rect 424 215 426 219
rect 365 208 367 213
rect 372 208 374 213
rect 332 206 357 208
rect 437 212 439 217
rect 444 212 446 217
rect 464 212 466 217
rect 471 212 473 217
rect 484 215 486 219
rect 504 215 506 219
rect 554 228 563 230
rect 579 230 581 233
rect 561 225 563 228
rect 571 225 573 229
rect 579 228 583 230
rect 581 225 583 228
rect 588 225 590 234
rect 629 233 635 235
rect 639 237 645 239
rect 639 235 641 237
rect 643 235 645 237
rect 639 233 645 235
rect 629 228 631 233
rect 642 228 644 233
rect 649 228 651 241
rect 669 228 671 241
rect 679 239 681 250
rect 689 239 691 243
rect 675 237 681 239
rect 675 235 677 237
rect 679 235 681 237
rect 675 233 681 235
rect 685 237 691 239
rect 685 235 687 237
rect 689 235 691 237
rect 685 233 691 235
rect 676 228 678 233
rect 689 228 691 233
rect 709 239 711 243
rect 719 239 721 250
rect 729 247 731 250
rect 729 245 735 247
rect 729 243 731 245
rect 733 243 735 245
rect 729 241 735 243
rect 743 245 749 247
rect 743 243 745 245
rect 747 243 749 245
rect 794 270 796 274
rect 774 261 776 265
rect 784 261 786 265
rect 848 261 850 265
rect 858 263 860 268
rect 868 263 870 268
rect 888 263 890 268
rect 898 263 900 268
rect 977 270 979 274
rect 908 261 910 265
rect 928 261 930 265
rect 938 263 940 268
rect 948 263 950 268
rect 743 241 749 243
rect 709 237 715 239
rect 709 235 711 237
rect 713 235 715 237
rect 709 233 715 235
rect 719 237 725 239
rect 719 235 721 237
rect 723 235 725 237
rect 719 233 725 235
rect 709 228 711 233
rect 722 228 724 233
rect 729 228 731 241
rect 747 240 749 241
rect 758 240 760 243
rect 774 240 776 243
rect 747 238 760 240
rect 766 238 776 240
rect 784 239 786 243
rect 794 240 796 243
rect 750 230 752 238
rect 766 234 768 238
rect 759 232 768 234
rect 780 237 786 239
rect 780 235 782 237
rect 784 235 786 237
rect 780 233 786 235
rect 790 238 796 240
rect 790 236 792 238
rect 794 236 796 238
rect 790 234 796 236
rect 848 239 850 243
rect 858 239 860 250
rect 868 247 870 250
rect 888 247 890 250
rect 868 245 874 247
rect 868 243 870 245
rect 872 243 874 245
rect 868 241 874 243
rect 884 245 890 247
rect 884 243 886 245
rect 888 243 890 245
rect 884 241 890 243
rect 848 237 854 239
rect 848 235 850 237
rect 852 235 854 237
rect 759 230 761 232
rect 763 230 768 232
rect 545 218 547 221
rect 517 212 519 217
rect 524 212 526 217
rect 545 216 550 218
rect 548 208 550 216
rect 561 212 563 216
rect 571 208 573 216
rect 629 215 631 219
rect 581 208 583 213
rect 588 208 590 213
rect 548 206 573 208
rect 642 212 644 217
rect 649 212 651 217
rect 669 212 671 217
rect 676 212 678 217
rect 689 215 691 219
rect 709 215 711 219
rect 759 228 768 230
rect 784 230 786 233
rect 766 225 768 228
rect 776 225 778 229
rect 784 228 788 230
rect 786 225 788 228
rect 793 225 795 234
rect 848 233 854 235
rect 858 237 864 239
rect 858 235 860 237
rect 862 235 864 237
rect 858 233 864 235
rect 848 228 850 233
rect 861 228 863 233
rect 868 228 870 241
rect 888 228 890 241
rect 898 239 900 250
rect 908 239 910 243
rect 894 237 900 239
rect 894 235 896 237
rect 898 235 900 237
rect 894 233 900 235
rect 904 237 910 239
rect 904 235 906 237
rect 908 235 910 237
rect 904 233 910 235
rect 895 228 897 233
rect 908 228 910 233
rect 928 239 930 243
rect 938 239 940 250
rect 948 247 950 250
rect 948 245 954 247
rect 948 243 950 245
rect 952 243 954 245
rect 948 241 954 243
rect 962 245 968 247
rect 962 243 964 245
rect 966 243 968 245
rect 1013 270 1015 274
rect 993 261 995 265
rect 1003 261 1005 265
rect 1101 270 1103 274
rect 1052 261 1054 265
rect 1062 263 1064 268
rect 1072 263 1074 268
rect 962 241 968 243
rect 928 237 934 239
rect 928 235 930 237
rect 932 235 934 237
rect 928 233 934 235
rect 938 237 944 239
rect 938 235 940 237
rect 942 235 944 237
rect 938 233 944 235
rect 928 228 930 233
rect 941 228 943 233
rect 948 228 950 241
rect 966 240 968 241
rect 977 240 979 243
rect 993 240 995 243
rect 966 238 979 240
rect 985 238 995 240
rect 1003 239 1005 243
rect 1013 240 1015 243
rect 969 230 971 238
rect 985 234 987 238
rect 978 232 987 234
rect 999 237 1005 239
rect 999 235 1001 237
rect 1003 235 1005 237
rect 999 233 1005 235
rect 1009 238 1015 240
rect 1009 236 1011 238
rect 1013 236 1015 238
rect 1009 234 1015 236
rect 1052 239 1054 243
rect 1062 239 1064 250
rect 1072 247 1074 250
rect 1072 245 1078 247
rect 1072 243 1074 245
rect 1076 243 1078 245
rect 1072 241 1078 243
rect 1086 245 1092 247
rect 1086 243 1088 245
rect 1090 243 1092 245
rect 1137 270 1139 274
rect 1117 261 1119 265
rect 1127 261 1129 265
rect 1086 241 1092 243
rect 1052 237 1058 239
rect 1052 235 1054 237
rect 1056 235 1058 237
rect 978 230 980 232
rect 982 230 987 232
rect 750 218 752 221
rect 722 212 724 217
rect 729 212 731 217
rect 750 216 755 218
rect 753 208 755 216
rect 766 212 768 216
rect 776 208 778 216
rect 848 215 850 219
rect 786 208 788 213
rect 793 208 795 213
rect 753 206 778 208
rect 861 212 863 217
rect 868 212 870 217
rect 888 212 890 217
rect 895 212 897 217
rect 908 215 910 219
rect 928 215 930 219
rect 978 228 987 230
rect 1003 230 1005 233
rect 985 225 987 228
rect 995 225 997 229
rect 1003 228 1007 230
rect 1005 225 1007 228
rect 1012 225 1014 234
rect 1052 233 1058 235
rect 1062 237 1068 239
rect 1062 235 1064 237
rect 1066 235 1068 237
rect 1062 233 1068 235
rect 1052 228 1054 233
rect 1065 228 1067 233
rect 1072 228 1074 241
rect 1090 240 1092 241
rect 1101 240 1103 243
rect 1117 240 1119 243
rect 1090 238 1103 240
rect 1109 238 1119 240
rect 1127 239 1129 243
rect 1137 240 1139 243
rect 1093 230 1095 238
rect 1109 234 1111 238
rect 1102 232 1111 234
rect 1123 237 1129 239
rect 1123 235 1125 237
rect 1127 235 1129 237
rect 1123 233 1129 235
rect 1133 238 1139 240
rect 1133 236 1135 238
rect 1137 236 1139 238
rect 1133 234 1139 236
rect 1102 230 1104 232
rect 1106 230 1111 232
rect 969 218 971 221
rect 941 212 943 217
rect 948 212 950 217
rect 969 216 974 218
rect 972 208 974 216
rect 985 212 987 216
rect 995 208 997 216
rect 1052 215 1054 219
rect 1102 228 1111 230
rect 1127 230 1129 233
rect 1109 225 1111 228
rect 1119 225 1121 229
rect 1127 228 1131 230
rect 1129 225 1131 228
rect 1136 225 1138 234
rect 1093 218 1095 221
rect 1005 208 1007 213
rect 1012 208 1014 213
rect 972 206 997 208
rect 1065 212 1067 217
rect 1072 212 1074 217
rect 1093 216 1098 218
rect 1096 208 1098 216
rect 1109 212 1111 216
rect 1119 208 1121 216
rect 1129 208 1131 213
rect 1136 208 1138 213
rect 1096 206 1121 208
rect 158 187 160 192
rect 168 184 170 189
rect 178 184 180 189
rect 198 189 200 193
rect 211 191 213 196
rect 218 191 220 196
rect 242 200 267 202
rect 242 192 244 200
rect 255 192 257 196
rect 265 192 267 200
rect 275 195 277 200
rect 282 195 284 200
rect 239 190 244 192
rect 239 187 241 190
rect 158 175 160 178
rect 168 175 170 178
rect 158 173 164 175
rect 158 171 160 173
rect 162 171 164 173
rect 158 169 164 171
rect 168 173 174 175
rect 168 171 170 173
rect 172 171 174 173
rect 168 169 174 171
rect 158 166 160 169
rect 171 159 173 169
rect 178 168 180 178
rect 198 175 200 180
rect 211 175 213 180
rect 198 173 204 175
rect 198 171 200 173
rect 202 171 204 173
rect 198 169 204 171
rect 208 173 214 175
rect 208 171 210 173
rect 212 171 214 173
rect 208 169 214 171
rect 178 166 184 168
rect 178 164 180 166
rect 182 164 184 166
rect 198 165 200 169
rect 178 162 184 164
rect 178 159 180 162
rect 158 143 160 148
rect 208 158 210 169
rect 218 167 220 180
rect 303 189 305 193
rect 316 191 318 196
rect 323 191 325 196
rect 347 200 372 202
rect 347 192 349 200
rect 360 192 362 196
rect 370 192 372 200
rect 380 195 382 200
rect 387 195 389 200
rect 255 180 257 183
rect 248 178 257 180
rect 265 179 267 183
rect 275 180 277 183
rect 239 170 241 178
rect 248 176 250 178
rect 252 176 257 178
rect 248 174 257 176
rect 273 178 277 180
rect 273 175 275 178
rect 255 170 257 174
rect 269 173 275 175
rect 282 174 284 183
rect 344 190 349 192
rect 344 187 346 190
rect 303 175 305 180
rect 316 175 318 180
rect 269 171 271 173
rect 273 171 275 173
rect 236 168 249 170
rect 255 168 265 170
rect 269 169 275 171
rect 236 167 238 168
rect 218 165 224 167
rect 218 163 220 165
rect 222 163 224 165
rect 218 161 224 163
rect 232 165 238 167
rect 247 165 249 168
rect 263 165 265 168
rect 273 165 275 169
rect 279 172 285 174
rect 279 170 281 172
rect 283 170 285 172
rect 279 168 285 170
rect 283 165 285 168
rect 303 173 309 175
rect 303 171 305 173
rect 307 171 309 173
rect 303 169 309 171
rect 313 173 319 175
rect 313 171 315 173
rect 317 171 319 173
rect 313 169 319 171
rect 303 165 305 169
rect 232 163 234 165
rect 236 163 238 165
rect 232 161 238 163
rect 218 158 220 161
rect 198 143 200 147
rect 208 140 210 145
rect 218 140 220 145
rect 171 134 173 138
rect 178 134 180 138
rect 263 143 265 147
rect 273 143 275 147
rect 247 134 249 138
rect 313 158 315 169
rect 323 167 325 180
rect 408 187 410 192
rect 360 180 362 183
rect 353 178 362 180
rect 370 179 372 183
rect 380 180 382 183
rect 344 170 346 178
rect 353 176 355 178
rect 357 176 362 178
rect 353 174 362 176
rect 378 178 382 180
rect 378 175 380 178
rect 360 170 362 174
rect 374 173 380 175
rect 387 174 389 183
rect 418 184 420 189
rect 428 184 430 189
rect 448 189 450 193
rect 461 191 463 196
rect 468 191 470 196
rect 492 200 517 202
rect 492 192 494 200
rect 505 192 507 196
rect 515 192 517 200
rect 525 195 527 200
rect 532 195 534 200
rect 489 190 494 192
rect 489 187 491 190
rect 408 175 410 178
rect 418 175 420 178
rect 374 171 376 173
rect 378 171 380 173
rect 341 168 354 170
rect 360 168 370 170
rect 374 169 380 171
rect 341 167 343 168
rect 323 165 329 167
rect 323 163 325 165
rect 327 163 329 165
rect 323 161 329 163
rect 337 165 343 167
rect 352 165 354 168
rect 368 165 370 168
rect 378 165 380 169
rect 384 172 390 174
rect 384 170 386 172
rect 388 170 390 172
rect 384 168 390 170
rect 388 165 390 168
rect 408 173 414 175
rect 408 171 410 173
rect 412 171 414 173
rect 408 169 414 171
rect 418 173 424 175
rect 418 171 420 173
rect 422 171 424 173
rect 418 169 424 171
rect 408 166 410 169
rect 337 163 339 165
rect 341 163 343 165
rect 337 161 343 163
rect 323 158 325 161
rect 303 143 305 147
rect 313 140 315 145
rect 323 140 325 145
rect 283 134 285 138
rect 368 143 370 147
rect 378 143 380 147
rect 352 134 354 138
rect 421 159 423 169
rect 428 168 430 178
rect 448 175 450 180
rect 461 175 463 180
rect 448 173 454 175
rect 448 171 450 173
rect 452 171 454 173
rect 448 169 454 171
rect 458 173 464 175
rect 458 171 460 173
rect 462 171 464 173
rect 458 169 464 171
rect 428 166 434 168
rect 428 164 430 166
rect 432 164 434 166
rect 448 165 450 169
rect 428 162 434 164
rect 428 159 430 162
rect 408 143 410 148
rect 388 134 390 138
rect 458 158 460 169
rect 468 167 470 180
rect 553 189 555 193
rect 566 191 568 196
rect 573 191 575 196
rect 597 200 622 202
rect 597 192 599 200
rect 610 192 612 196
rect 620 192 622 200
rect 630 195 632 200
rect 637 195 639 200
rect 505 180 507 183
rect 498 178 507 180
rect 515 179 517 183
rect 525 180 527 183
rect 489 170 491 178
rect 498 176 500 178
rect 502 176 507 178
rect 498 174 507 176
rect 523 178 527 180
rect 523 175 525 178
rect 505 170 507 174
rect 519 173 525 175
rect 532 174 534 183
rect 594 190 599 192
rect 594 187 596 190
rect 553 175 555 180
rect 566 175 568 180
rect 519 171 521 173
rect 523 171 525 173
rect 486 168 499 170
rect 505 168 515 170
rect 519 169 525 171
rect 486 167 488 168
rect 468 165 474 167
rect 468 163 470 165
rect 472 163 474 165
rect 468 161 474 163
rect 482 165 488 167
rect 497 165 499 168
rect 513 165 515 168
rect 523 165 525 169
rect 529 172 535 174
rect 529 170 531 172
rect 533 170 535 172
rect 529 168 535 170
rect 533 165 535 168
rect 553 173 559 175
rect 553 171 555 173
rect 557 171 559 173
rect 553 169 559 171
rect 563 173 569 175
rect 563 171 565 173
rect 567 171 569 173
rect 563 169 569 171
rect 553 165 555 169
rect 482 163 484 165
rect 486 163 488 165
rect 482 161 488 163
rect 468 158 470 161
rect 448 143 450 147
rect 458 140 460 145
rect 468 140 470 145
rect 421 134 423 138
rect 428 134 430 138
rect 513 143 515 147
rect 523 143 525 147
rect 497 134 499 138
rect 563 158 565 169
rect 573 167 575 180
rect 658 187 660 192
rect 610 180 612 183
rect 603 178 612 180
rect 620 179 622 183
rect 630 180 632 183
rect 594 170 596 178
rect 603 176 605 178
rect 607 176 612 178
rect 603 174 612 176
rect 628 178 632 180
rect 628 175 630 178
rect 610 170 612 174
rect 624 173 630 175
rect 637 174 639 183
rect 668 184 670 189
rect 678 184 680 189
rect 698 189 700 193
rect 711 191 713 196
rect 718 191 720 196
rect 742 200 767 202
rect 742 192 744 200
rect 755 192 757 196
rect 765 192 767 200
rect 775 195 777 200
rect 782 195 784 200
rect 739 190 744 192
rect 739 187 741 190
rect 658 175 660 178
rect 668 175 670 178
rect 624 171 626 173
rect 628 171 630 173
rect 591 168 604 170
rect 610 168 620 170
rect 624 169 630 171
rect 591 167 593 168
rect 573 165 579 167
rect 573 163 575 165
rect 577 163 579 165
rect 573 161 579 163
rect 587 165 593 167
rect 602 165 604 168
rect 618 165 620 168
rect 628 165 630 169
rect 634 172 640 174
rect 634 170 636 172
rect 638 170 640 172
rect 634 168 640 170
rect 638 165 640 168
rect 658 173 664 175
rect 658 171 660 173
rect 662 171 664 173
rect 658 169 664 171
rect 668 173 674 175
rect 668 171 670 173
rect 672 171 674 173
rect 668 169 674 171
rect 658 166 660 169
rect 587 163 589 165
rect 591 163 593 165
rect 587 161 593 163
rect 573 158 575 161
rect 553 143 555 147
rect 563 140 565 145
rect 573 140 575 145
rect 533 134 535 138
rect 618 143 620 147
rect 628 143 630 147
rect 602 134 604 138
rect 671 159 673 169
rect 678 168 680 178
rect 698 175 700 180
rect 711 175 713 180
rect 698 173 704 175
rect 698 171 700 173
rect 702 171 704 173
rect 698 169 704 171
rect 708 173 714 175
rect 708 171 710 173
rect 712 171 714 173
rect 708 169 714 171
rect 678 166 684 168
rect 678 164 680 166
rect 682 164 684 166
rect 698 165 700 169
rect 678 162 684 164
rect 678 159 680 162
rect 658 143 660 148
rect 638 134 640 138
rect 708 158 710 169
rect 718 167 720 180
rect 803 189 805 193
rect 816 191 818 196
rect 823 191 825 196
rect 847 200 872 202
rect 847 192 849 200
rect 860 192 862 196
rect 870 192 872 200
rect 880 195 882 200
rect 887 195 889 200
rect 755 180 757 183
rect 748 178 757 180
rect 765 179 767 183
rect 775 180 777 183
rect 739 170 741 178
rect 748 176 750 178
rect 752 176 757 178
rect 748 174 757 176
rect 773 178 777 180
rect 773 175 775 178
rect 755 170 757 174
rect 769 173 775 175
rect 782 174 784 183
rect 844 190 849 192
rect 844 187 846 190
rect 803 175 805 180
rect 816 175 818 180
rect 769 171 771 173
rect 773 171 775 173
rect 736 168 749 170
rect 755 168 765 170
rect 769 169 775 171
rect 736 167 738 168
rect 718 165 724 167
rect 718 163 720 165
rect 722 163 724 165
rect 718 161 724 163
rect 732 165 738 167
rect 747 165 749 168
rect 763 165 765 168
rect 773 165 775 169
rect 779 172 785 174
rect 779 170 781 172
rect 783 170 785 172
rect 779 168 785 170
rect 783 165 785 168
rect 803 173 809 175
rect 803 171 805 173
rect 807 171 809 173
rect 803 169 809 171
rect 813 173 819 175
rect 813 171 815 173
rect 817 171 819 173
rect 813 169 819 171
rect 803 165 805 169
rect 732 163 734 165
rect 736 163 738 165
rect 732 161 738 163
rect 718 158 720 161
rect 698 143 700 147
rect 708 140 710 145
rect 718 140 720 145
rect 671 134 673 138
rect 678 134 680 138
rect 763 143 765 147
rect 773 143 775 147
rect 747 134 749 138
rect 813 158 815 169
rect 823 167 825 180
rect 908 187 910 192
rect 860 180 862 183
rect 853 178 862 180
rect 870 179 872 183
rect 880 180 882 183
rect 844 170 846 178
rect 853 176 855 178
rect 857 176 862 178
rect 853 174 862 176
rect 878 178 882 180
rect 878 175 880 178
rect 860 170 862 174
rect 874 173 880 175
rect 887 174 889 183
rect 918 184 920 189
rect 928 184 930 189
rect 948 189 950 193
rect 961 191 963 196
rect 968 191 970 196
rect 992 200 1017 202
rect 992 192 994 200
rect 1005 192 1007 196
rect 1015 192 1017 200
rect 1025 195 1027 200
rect 1032 195 1034 200
rect 989 190 994 192
rect 989 187 991 190
rect 908 175 910 178
rect 918 175 920 178
rect 874 171 876 173
rect 878 171 880 173
rect 841 168 854 170
rect 860 168 870 170
rect 874 169 880 171
rect 841 167 843 168
rect 823 165 829 167
rect 823 163 825 165
rect 827 163 829 165
rect 823 161 829 163
rect 837 165 843 167
rect 852 165 854 168
rect 868 165 870 168
rect 878 165 880 169
rect 884 172 890 174
rect 884 170 886 172
rect 888 170 890 172
rect 884 168 890 170
rect 888 165 890 168
rect 908 173 914 175
rect 908 171 910 173
rect 912 171 914 173
rect 908 169 914 171
rect 918 173 924 175
rect 918 171 920 173
rect 922 171 924 173
rect 918 169 924 171
rect 908 166 910 169
rect 837 163 839 165
rect 841 163 843 165
rect 837 161 843 163
rect 823 158 825 161
rect 803 143 805 147
rect 813 140 815 145
rect 823 140 825 145
rect 783 134 785 138
rect 868 143 870 147
rect 878 143 880 147
rect 852 134 854 138
rect 921 159 923 169
rect 928 168 930 178
rect 948 175 950 180
rect 961 175 963 180
rect 948 173 954 175
rect 948 171 950 173
rect 952 171 954 173
rect 948 169 954 171
rect 958 173 964 175
rect 958 171 960 173
rect 962 171 964 173
rect 958 169 964 171
rect 928 166 934 168
rect 928 164 930 166
rect 932 164 934 166
rect 948 165 950 169
rect 928 162 934 164
rect 928 159 930 162
rect 908 143 910 148
rect 888 134 890 138
rect 958 158 960 169
rect 968 167 970 180
rect 1053 189 1055 193
rect 1066 191 1068 196
rect 1073 191 1075 196
rect 1097 200 1122 202
rect 1097 192 1099 200
rect 1110 192 1112 196
rect 1120 192 1122 200
rect 1130 195 1132 200
rect 1137 195 1139 200
rect 1005 180 1007 183
rect 998 178 1007 180
rect 1015 179 1017 183
rect 1025 180 1027 183
rect 989 170 991 178
rect 998 176 1000 178
rect 1002 176 1007 178
rect 998 174 1007 176
rect 1023 178 1027 180
rect 1023 175 1025 178
rect 1005 170 1007 174
rect 1019 173 1025 175
rect 1032 174 1034 183
rect 1094 190 1099 192
rect 1094 187 1096 190
rect 1053 175 1055 180
rect 1066 175 1068 180
rect 1019 171 1021 173
rect 1023 171 1025 173
rect 986 168 999 170
rect 1005 168 1015 170
rect 1019 169 1025 171
rect 986 167 988 168
rect 968 165 974 167
rect 968 163 970 165
rect 972 163 974 165
rect 968 161 974 163
rect 982 165 988 167
rect 997 165 999 168
rect 1013 165 1015 168
rect 1023 165 1025 169
rect 1029 172 1035 174
rect 1029 170 1031 172
rect 1033 170 1035 172
rect 1029 168 1035 170
rect 1033 165 1035 168
rect 1053 173 1059 175
rect 1053 171 1055 173
rect 1057 171 1059 173
rect 1053 169 1059 171
rect 1063 173 1069 175
rect 1063 171 1065 173
rect 1067 171 1069 173
rect 1063 169 1069 171
rect 1053 165 1055 169
rect 982 163 984 165
rect 986 163 988 165
rect 982 161 988 163
rect 968 158 970 161
rect 948 143 950 147
rect 958 140 960 145
rect 968 140 970 145
rect 921 134 923 138
rect 928 134 930 138
rect 1013 143 1015 147
rect 1023 143 1025 147
rect 997 134 999 138
rect 1063 158 1065 169
rect 1073 167 1075 180
rect 1110 180 1112 183
rect 1103 178 1112 180
rect 1120 179 1122 183
rect 1130 180 1132 183
rect 1094 170 1096 178
rect 1103 176 1105 178
rect 1107 176 1112 178
rect 1103 174 1112 176
rect 1128 178 1132 180
rect 1128 175 1130 178
rect 1110 170 1112 174
rect 1124 173 1130 175
rect 1137 174 1139 183
rect 1124 171 1126 173
rect 1128 171 1130 173
rect 1091 168 1104 170
rect 1110 168 1120 170
rect 1124 169 1130 171
rect 1091 167 1093 168
rect 1073 165 1079 167
rect 1073 163 1075 165
rect 1077 163 1079 165
rect 1073 161 1079 163
rect 1087 165 1093 167
rect 1102 165 1104 168
rect 1118 165 1120 168
rect 1128 165 1130 169
rect 1134 172 1140 174
rect 1134 170 1136 172
rect 1138 170 1140 172
rect 1134 168 1140 170
rect 1138 165 1140 168
rect 1087 163 1089 165
rect 1091 163 1093 165
rect 1087 161 1093 163
rect 1073 158 1075 161
rect 1053 143 1055 147
rect 1063 140 1065 145
rect 1073 140 1075 145
rect 1033 134 1035 138
rect 1118 143 1120 147
rect 1128 143 1130 147
rect 1102 134 1104 138
rect 1138 134 1140 138
rect 170 126 172 130
rect 177 126 179 130
rect 157 116 159 121
rect 246 126 248 130
rect 197 117 199 121
rect 207 119 209 124
rect 217 119 219 124
rect 157 95 159 98
rect 170 95 172 105
rect 177 102 179 105
rect 177 100 183 102
rect 177 98 179 100
rect 181 98 183 100
rect 177 96 183 98
rect 157 93 163 95
rect 157 91 159 93
rect 161 91 163 93
rect 157 89 163 91
rect 167 93 173 95
rect 167 91 169 93
rect 171 91 173 93
rect 167 89 173 91
rect 157 86 159 89
rect 167 86 169 89
rect 177 86 179 96
rect 197 95 199 99
rect 207 95 209 106
rect 217 103 219 106
rect 217 101 223 103
rect 217 99 219 101
rect 221 99 223 101
rect 217 97 223 99
rect 231 101 237 103
rect 231 99 233 101
rect 235 99 237 101
rect 282 126 284 130
rect 262 117 264 121
rect 272 117 274 121
rect 351 126 353 130
rect 302 117 304 121
rect 312 119 314 124
rect 322 119 324 124
rect 231 97 237 99
rect 197 93 203 95
rect 197 91 199 93
rect 201 91 203 93
rect 197 89 203 91
rect 207 93 213 95
rect 207 91 209 93
rect 211 91 213 93
rect 207 89 213 91
rect 197 84 199 89
rect 210 84 212 89
rect 217 84 219 97
rect 235 96 237 97
rect 246 96 248 99
rect 262 96 264 99
rect 235 94 248 96
rect 254 94 264 96
rect 272 95 274 99
rect 282 96 284 99
rect 238 86 240 94
rect 254 90 256 94
rect 247 88 256 90
rect 268 93 274 95
rect 268 91 270 93
rect 272 91 274 93
rect 268 89 274 91
rect 278 94 284 96
rect 278 92 280 94
rect 282 92 284 94
rect 278 90 284 92
rect 302 95 304 99
rect 312 95 314 106
rect 322 103 324 106
rect 322 101 328 103
rect 322 99 324 101
rect 326 99 328 101
rect 322 97 328 99
rect 336 101 342 103
rect 336 99 338 101
rect 340 99 342 101
rect 387 126 389 130
rect 367 117 369 121
rect 377 117 379 121
rect 420 126 422 130
rect 427 126 429 130
rect 407 116 409 121
rect 336 97 342 99
rect 302 93 308 95
rect 302 91 304 93
rect 306 91 308 93
rect 247 86 249 88
rect 251 86 256 88
rect 157 72 159 77
rect 167 75 169 80
rect 177 75 179 80
rect 197 71 199 75
rect 247 84 256 86
rect 272 86 274 89
rect 254 81 256 84
rect 264 81 266 85
rect 272 84 276 86
rect 274 81 276 84
rect 281 81 283 90
rect 302 89 308 91
rect 312 93 318 95
rect 312 91 314 93
rect 316 91 318 93
rect 312 89 318 91
rect 302 84 304 89
rect 315 84 317 89
rect 322 84 324 97
rect 340 96 342 97
rect 351 96 353 99
rect 367 96 369 99
rect 340 94 353 96
rect 359 94 369 96
rect 377 95 379 99
rect 387 96 389 99
rect 496 126 498 130
rect 447 117 449 121
rect 457 119 459 124
rect 467 119 469 124
rect 343 86 345 94
rect 359 90 361 94
rect 352 88 361 90
rect 373 93 379 95
rect 373 91 375 93
rect 377 91 379 93
rect 373 89 379 91
rect 383 94 389 96
rect 383 92 385 94
rect 387 92 389 94
rect 383 90 389 92
rect 407 95 409 98
rect 420 95 422 105
rect 427 102 429 105
rect 427 100 433 102
rect 427 98 429 100
rect 431 98 433 100
rect 427 96 433 98
rect 407 93 413 95
rect 407 91 409 93
rect 411 91 413 93
rect 352 86 354 88
rect 356 86 361 88
rect 238 74 240 77
rect 210 68 212 73
rect 217 68 219 73
rect 238 72 243 74
rect 241 64 243 72
rect 254 68 256 72
rect 264 64 266 72
rect 302 71 304 75
rect 352 84 361 86
rect 377 86 379 89
rect 359 81 361 84
rect 369 81 371 85
rect 377 84 381 86
rect 379 81 381 84
rect 386 81 388 90
rect 407 89 413 91
rect 417 93 423 95
rect 417 91 419 93
rect 421 91 423 93
rect 417 89 423 91
rect 407 86 409 89
rect 417 86 419 89
rect 427 86 429 96
rect 447 95 449 99
rect 457 95 459 106
rect 467 103 469 106
rect 467 101 473 103
rect 467 99 469 101
rect 471 99 473 101
rect 467 97 473 99
rect 481 101 487 103
rect 481 99 483 101
rect 485 99 487 101
rect 532 126 534 130
rect 512 117 514 121
rect 522 117 524 121
rect 601 126 603 130
rect 552 117 554 121
rect 562 119 564 124
rect 572 119 574 124
rect 481 97 487 99
rect 447 93 453 95
rect 447 91 449 93
rect 451 91 453 93
rect 447 89 453 91
rect 457 93 463 95
rect 457 91 459 93
rect 461 91 463 93
rect 457 89 463 91
rect 343 74 345 77
rect 274 64 276 69
rect 281 64 283 69
rect 241 62 266 64
rect 315 68 317 73
rect 322 68 324 73
rect 343 72 348 74
rect 346 64 348 72
rect 359 68 361 72
rect 369 64 371 72
rect 447 84 449 89
rect 460 84 462 89
rect 467 84 469 97
rect 485 96 487 97
rect 496 96 498 99
rect 512 96 514 99
rect 485 94 498 96
rect 504 94 514 96
rect 522 95 524 99
rect 532 96 534 99
rect 488 86 490 94
rect 504 90 506 94
rect 497 88 506 90
rect 518 93 524 95
rect 518 91 520 93
rect 522 91 524 93
rect 518 89 524 91
rect 528 94 534 96
rect 528 92 530 94
rect 532 92 534 94
rect 528 90 534 92
rect 552 95 554 99
rect 562 95 564 106
rect 572 103 574 106
rect 572 101 578 103
rect 572 99 574 101
rect 576 99 578 101
rect 572 97 578 99
rect 586 101 592 103
rect 586 99 588 101
rect 590 99 592 101
rect 637 126 639 130
rect 617 117 619 121
rect 627 117 629 121
rect 670 126 672 130
rect 677 126 679 130
rect 657 116 659 121
rect 586 97 592 99
rect 552 93 558 95
rect 552 91 554 93
rect 556 91 558 93
rect 497 86 499 88
rect 501 86 506 88
rect 407 72 409 77
rect 417 75 419 80
rect 427 75 429 80
rect 379 64 381 69
rect 386 64 388 69
rect 346 62 371 64
rect 447 71 449 75
rect 497 84 506 86
rect 522 86 524 89
rect 504 81 506 84
rect 514 81 516 85
rect 522 84 526 86
rect 524 81 526 84
rect 531 81 533 90
rect 552 89 558 91
rect 562 93 568 95
rect 562 91 564 93
rect 566 91 568 93
rect 562 89 568 91
rect 552 84 554 89
rect 565 84 567 89
rect 572 84 574 97
rect 590 96 592 97
rect 601 96 603 99
rect 617 96 619 99
rect 590 94 603 96
rect 609 94 619 96
rect 627 95 629 99
rect 637 96 639 99
rect 746 126 748 130
rect 697 117 699 121
rect 707 119 709 124
rect 717 119 719 124
rect 593 86 595 94
rect 609 90 611 94
rect 602 88 611 90
rect 623 93 629 95
rect 623 91 625 93
rect 627 91 629 93
rect 623 89 629 91
rect 633 94 639 96
rect 633 92 635 94
rect 637 92 639 94
rect 633 90 639 92
rect 657 95 659 98
rect 670 95 672 105
rect 677 102 679 105
rect 677 100 683 102
rect 677 98 679 100
rect 681 98 683 100
rect 677 96 683 98
rect 657 93 663 95
rect 657 91 659 93
rect 661 91 663 93
rect 602 86 604 88
rect 606 86 611 88
rect 488 74 490 77
rect 460 68 462 73
rect 467 68 469 73
rect 488 72 493 74
rect 491 64 493 72
rect 504 68 506 72
rect 514 64 516 72
rect 552 71 554 75
rect 602 84 611 86
rect 627 86 629 89
rect 609 81 611 84
rect 619 81 621 85
rect 627 84 631 86
rect 629 81 631 84
rect 636 81 638 90
rect 657 89 663 91
rect 667 93 673 95
rect 667 91 669 93
rect 671 91 673 93
rect 667 89 673 91
rect 657 86 659 89
rect 667 86 669 89
rect 677 86 679 96
rect 697 95 699 99
rect 707 95 709 106
rect 717 103 719 106
rect 717 101 723 103
rect 717 99 719 101
rect 721 99 723 101
rect 717 97 723 99
rect 731 101 737 103
rect 731 99 733 101
rect 735 99 737 101
rect 782 126 784 130
rect 762 117 764 121
rect 772 117 774 121
rect 851 126 853 130
rect 802 117 804 121
rect 812 119 814 124
rect 822 119 824 124
rect 731 97 737 99
rect 697 93 703 95
rect 697 91 699 93
rect 701 91 703 93
rect 697 89 703 91
rect 707 93 713 95
rect 707 91 709 93
rect 711 91 713 93
rect 707 89 713 91
rect 593 74 595 77
rect 524 64 526 69
rect 531 64 533 69
rect 491 62 516 64
rect 565 68 567 73
rect 572 68 574 73
rect 593 72 598 74
rect 596 64 598 72
rect 609 68 611 72
rect 619 64 621 72
rect 697 84 699 89
rect 710 84 712 89
rect 717 84 719 97
rect 735 96 737 97
rect 746 96 748 99
rect 762 96 764 99
rect 735 94 748 96
rect 754 94 764 96
rect 772 95 774 99
rect 782 96 784 99
rect 738 86 740 94
rect 754 90 756 94
rect 747 88 756 90
rect 768 93 774 95
rect 768 91 770 93
rect 772 91 774 93
rect 768 89 774 91
rect 778 94 784 96
rect 778 92 780 94
rect 782 92 784 94
rect 778 90 784 92
rect 802 95 804 99
rect 812 95 814 106
rect 822 103 824 106
rect 822 101 828 103
rect 822 99 824 101
rect 826 99 828 101
rect 822 97 828 99
rect 836 101 842 103
rect 836 99 838 101
rect 840 99 842 101
rect 887 126 889 130
rect 867 117 869 121
rect 877 117 879 121
rect 920 126 922 130
rect 927 126 929 130
rect 907 116 909 121
rect 836 97 842 99
rect 802 93 808 95
rect 802 91 804 93
rect 806 91 808 93
rect 747 86 749 88
rect 751 86 756 88
rect 657 72 659 77
rect 667 75 669 80
rect 677 75 679 80
rect 629 64 631 69
rect 636 64 638 69
rect 596 62 621 64
rect 697 71 699 75
rect 747 84 756 86
rect 772 86 774 89
rect 754 81 756 84
rect 764 81 766 85
rect 772 84 776 86
rect 774 81 776 84
rect 781 81 783 90
rect 802 89 808 91
rect 812 93 818 95
rect 812 91 814 93
rect 816 91 818 93
rect 812 89 818 91
rect 802 84 804 89
rect 815 84 817 89
rect 822 84 824 97
rect 840 96 842 97
rect 851 96 853 99
rect 867 96 869 99
rect 840 94 853 96
rect 859 94 869 96
rect 877 95 879 99
rect 887 96 889 99
rect 996 126 998 130
rect 947 117 949 121
rect 957 119 959 124
rect 967 119 969 124
rect 843 86 845 94
rect 859 90 861 94
rect 852 88 861 90
rect 873 93 879 95
rect 873 91 875 93
rect 877 91 879 93
rect 873 89 879 91
rect 883 94 889 96
rect 883 92 885 94
rect 887 92 889 94
rect 883 90 889 92
rect 907 95 909 98
rect 920 95 922 105
rect 927 102 929 105
rect 927 100 933 102
rect 927 98 929 100
rect 931 98 933 100
rect 927 96 933 98
rect 907 93 913 95
rect 907 91 909 93
rect 911 91 913 93
rect 852 86 854 88
rect 856 86 861 88
rect 738 74 740 77
rect 710 68 712 73
rect 717 68 719 73
rect 738 72 743 74
rect 741 64 743 72
rect 754 68 756 72
rect 764 64 766 72
rect 802 71 804 75
rect 852 84 861 86
rect 877 86 879 89
rect 859 81 861 84
rect 869 81 871 85
rect 877 84 881 86
rect 879 81 881 84
rect 886 81 888 90
rect 907 89 913 91
rect 917 93 923 95
rect 917 91 919 93
rect 921 91 923 93
rect 917 89 923 91
rect 907 86 909 89
rect 917 86 919 89
rect 927 86 929 96
rect 947 95 949 99
rect 957 95 959 106
rect 967 103 969 106
rect 967 101 973 103
rect 967 99 969 101
rect 971 99 973 101
rect 967 97 973 99
rect 981 101 987 103
rect 981 99 983 101
rect 985 99 987 101
rect 1032 126 1034 130
rect 1012 117 1014 121
rect 1022 117 1024 121
rect 1101 126 1103 130
rect 1052 117 1054 121
rect 1062 119 1064 124
rect 1072 119 1074 124
rect 981 97 987 99
rect 947 93 953 95
rect 947 91 949 93
rect 951 91 953 93
rect 947 89 953 91
rect 957 93 963 95
rect 957 91 959 93
rect 961 91 963 93
rect 957 89 963 91
rect 843 74 845 77
rect 774 64 776 69
rect 781 64 783 69
rect 741 62 766 64
rect 815 68 817 73
rect 822 68 824 73
rect 843 72 848 74
rect 846 64 848 72
rect 859 68 861 72
rect 869 64 871 72
rect 947 84 949 89
rect 960 84 962 89
rect 967 84 969 97
rect 985 96 987 97
rect 996 96 998 99
rect 1012 96 1014 99
rect 985 94 998 96
rect 1004 94 1014 96
rect 1022 95 1024 99
rect 1032 96 1034 99
rect 988 86 990 94
rect 1004 90 1006 94
rect 997 88 1006 90
rect 1018 93 1024 95
rect 1018 91 1020 93
rect 1022 91 1024 93
rect 1018 89 1024 91
rect 1028 94 1034 96
rect 1028 92 1030 94
rect 1032 92 1034 94
rect 1028 90 1034 92
rect 1052 95 1054 99
rect 1062 95 1064 106
rect 1072 103 1074 106
rect 1072 101 1078 103
rect 1072 99 1074 101
rect 1076 99 1078 101
rect 1072 97 1078 99
rect 1086 101 1092 103
rect 1086 99 1088 101
rect 1090 99 1092 101
rect 1137 126 1139 130
rect 1117 117 1119 121
rect 1127 117 1129 121
rect 1086 97 1092 99
rect 1052 93 1058 95
rect 1052 91 1054 93
rect 1056 91 1058 93
rect 997 86 999 88
rect 1001 86 1006 88
rect 907 72 909 77
rect 917 75 919 80
rect 927 75 929 80
rect 879 64 881 69
rect 886 64 888 69
rect 846 62 871 64
rect 947 71 949 75
rect 997 84 1006 86
rect 1022 86 1024 89
rect 1004 81 1006 84
rect 1014 81 1016 85
rect 1022 84 1026 86
rect 1024 81 1026 84
rect 1031 81 1033 90
rect 1052 89 1058 91
rect 1062 93 1068 95
rect 1062 91 1064 93
rect 1066 91 1068 93
rect 1062 89 1068 91
rect 1052 84 1054 89
rect 1065 84 1067 89
rect 1072 84 1074 97
rect 1090 96 1092 97
rect 1101 96 1103 99
rect 1117 96 1119 99
rect 1090 94 1103 96
rect 1109 94 1119 96
rect 1127 95 1129 99
rect 1137 96 1139 99
rect 1093 86 1095 94
rect 1109 90 1111 94
rect 1102 88 1111 90
rect 1123 93 1129 95
rect 1123 91 1125 93
rect 1127 91 1129 93
rect 1123 89 1129 91
rect 1133 94 1139 96
rect 1133 92 1135 94
rect 1137 92 1139 94
rect 1133 90 1139 92
rect 1102 86 1104 88
rect 1106 86 1111 88
rect 988 74 990 77
rect 960 68 962 73
rect 967 68 969 73
rect 988 72 993 74
rect 991 64 993 72
rect 1004 68 1006 72
rect 1014 64 1016 72
rect 1052 71 1054 75
rect 1102 84 1111 86
rect 1127 86 1129 89
rect 1109 81 1111 84
rect 1119 81 1121 85
rect 1127 84 1131 86
rect 1129 81 1131 84
rect 1136 81 1138 90
rect 1093 74 1095 77
rect 1024 64 1026 69
rect 1031 64 1033 69
rect 991 62 1016 64
rect 1065 68 1067 73
rect 1072 68 1074 73
rect 1093 72 1098 74
rect 1096 64 1098 72
rect 1109 68 1111 72
rect 1119 64 1121 72
rect 1129 64 1131 69
rect 1136 64 1138 69
rect 1096 62 1121 64
rect 156 43 158 48
rect 166 40 168 45
rect 176 40 178 45
rect 196 45 198 49
rect 209 47 211 52
rect 216 47 218 52
rect 240 56 265 58
rect 240 48 242 56
rect 253 48 255 52
rect 263 48 265 56
rect 273 51 275 56
rect 280 51 282 56
rect 237 46 242 48
rect 237 43 239 46
rect 156 31 158 34
rect 166 31 168 34
rect 156 29 162 31
rect 156 27 158 29
rect 160 27 162 29
rect 156 25 162 27
rect 166 29 172 31
rect 166 27 168 29
rect 170 27 172 29
rect 166 25 172 27
rect 156 22 158 25
rect 169 15 171 25
rect 176 24 178 34
rect 196 31 198 36
rect 209 31 211 36
rect 196 29 202 31
rect 196 27 198 29
rect 200 27 202 29
rect 196 25 202 27
rect 206 29 212 31
rect 206 27 208 29
rect 210 27 212 29
rect 206 25 212 27
rect 176 22 182 24
rect 176 20 178 22
rect 180 20 182 22
rect 196 21 198 25
rect 176 18 182 20
rect 176 15 178 18
rect 156 -1 158 4
rect 206 14 208 25
rect 216 23 218 36
rect 301 45 303 49
rect 314 47 316 52
rect 321 47 323 52
rect 345 56 370 58
rect 345 48 347 56
rect 358 48 360 52
rect 368 48 370 56
rect 378 51 380 56
rect 385 51 387 56
rect 253 36 255 39
rect 246 34 255 36
rect 263 35 265 39
rect 273 36 275 39
rect 237 26 239 34
rect 246 32 248 34
rect 250 32 255 34
rect 246 30 255 32
rect 271 34 275 36
rect 271 31 273 34
rect 253 26 255 30
rect 267 29 273 31
rect 280 30 282 39
rect 342 46 347 48
rect 342 43 344 46
rect 301 31 303 36
rect 314 31 316 36
rect 267 27 269 29
rect 271 27 273 29
rect 234 24 247 26
rect 253 24 263 26
rect 267 25 273 27
rect 234 23 236 24
rect 216 21 222 23
rect 216 19 218 21
rect 220 19 222 21
rect 216 17 222 19
rect 230 21 236 23
rect 245 21 247 24
rect 261 21 263 24
rect 271 21 273 25
rect 277 28 283 30
rect 277 26 279 28
rect 281 26 283 28
rect 277 24 283 26
rect 281 21 283 24
rect 301 29 307 31
rect 301 27 303 29
rect 305 27 307 29
rect 301 25 307 27
rect 311 29 317 31
rect 311 27 313 29
rect 315 27 317 29
rect 311 25 317 27
rect 301 21 303 25
rect 230 19 232 21
rect 234 19 236 21
rect 230 17 236 19
rect 216 14 218 17
rect 196 -1 198 3
rect 206 -4 208 1
rect 216 -4 218 1
rect 169 -10 171 -6
rect 176 -10 178 -6
rect 261 -1 263 3
rect 271 -1 273 3
rect 245 -10 247 -6
rect 311 14 313 25
rect 321 23 323 36
rect 406 43 408 48
rect 358 36 360 39
rect 351 34 360 36
rect 368 35 370 39
rect 378 36 380 39
rect 342 26 344 34
rect 351 32 353 34
rect 355 32 360 34
rect 351 30 360 32
rect 376 34 380 36
rect 376 31 378 34
rect 358 26 360 30
rect 372 29 378 31
rect 385 30 387 39
rect 416 40 418 45
rect 426 40 428 45
rect 446 45 448 49
rect 459 47 461 52
rect 466 47 468 52
rect 490 56 515 58
rect 490 48 492 56
rect 503 48 505 52
rect 513 48 515 56
rect 523 51 525 56
rect 530 51 532 56
rect 487 46 492 48
rect 487 43 489 46
rect 406 31 408 34
rect 416 31 418 34
rect 372 27 374 29
rect 376 27 378 29
rect 339 24 352 26
rect 358 24 368 26
rect 372 25 378 27
rect 339 23 341 24
rect 321 21 327 23
rect 321 19 323 21
rect 325 19 327 21
rect 321 17 327 19
rect 335 21 341 23
rect 350 21 352 24
rect 366 21 368 24
rect 376 21 378 25
rect 382 28 388 30
rect 382 26 384 28
rect 386 26 388 28
rect 382 24 388 26
rect 386 21 388 24
rect 406 29 412 31
rect 406 27 408 29
rect 410 27 412 29
rect 406 25 412 27
rect 416 29 422 31
rect 416 27 418 29
rect 420 27 422 29
rect 416 25 422 27
rect 406 22 408 25
rect 335 19 337 21
rect 339 19 341 21
rect 335 17 341 19
rect 321 14 323 17
rect 301 -1 303 3
rect 311 -4 313 1
rect 321 -4 323 1
rect 281 -10 283 -6
rect 366 -1 368 3
rect 376 -1 378 3
rect 350 -10 352 -6
rect 419 15 421 25
rect 426 24 428 34
rect 446 31 448 36
rect 459 31 461 36
rect 446 29 452 31
rect 446 27 448 29
rect 450 27 452 29
rect 446 25 452 27
rect 456 29 462 31
rect 456 27 458 29
rect 460 27 462 29
rect 456 25 462 27
rect 426 22 432 24
rect 426 20 428 22
rect 430 20 432 22
rect 446 21 448 25
rect 426 18 432 20
rect 426 15 428 18
rect 406 -1 408 4
rect 386 -10 388 -6
rect 456 14 458 25
rect 466 23 468 36
rect 551 45 553 49
rect 564 47 566 52
rect 571 47 573 52
rect 595 56 620 58
rect 595 48 597 56
rect 608 48 610 52
rect 618 48 620 56
rect 628 51 630 56
rect 635 51 637 56
rect 503 36 505 39
rect 496 34 505 36
rect 513 35 515 39
rect 523 36 525 39
rect 487 26 489 34
rect 496 32 498 34
rect 500 32 505 34
rect 496 30 505 32
rect 521 34 525 36
rect 521 31 523 34
rect 503 26 505 30
rect 517 29 523 31
rect 530 30 532 39
rect 592 46 597 48
rect 592 43 594 46
rect 551 31 553 36
rect 564 31 566 36
rect 517 27 519 29
rect 521 27 523 29
rect 484 24 497 26
rect 503 24 513 26
rect 517 25 523 27
rect 484 23 486 24
rect 466 21 472 23
rect 466 19 468 21
rect 470 19 472 21
rect 466 17 472 19
rect 480 21 486 23
rect 495 21 497 24
rect 511 21 513 24
rect 521 21 523 25
rect 527 28 533 30
rect 527 26 529 28
rect 531 26 533 28
rect 527 24 533 26
rect 531 21 533 24
rect 551 29 557 31
rect 551 27 553 29
rect 555 27 557 29
rect 551 25 557 27
rect 561 29 567 31
rect 561 27 563 29
rect 565 27 567 29
rect 561 25 567 27
rect 551 21 553 25
rect 480 19 482 21
rect 484 19 486 21
rect 480 17 486 19
rect 466 14 468 17
rect 446 -1 448 3
rect 456 -4 458 1
rect 466 -4 468 1
rect 419 -10 421 -6
rect 426 -10 428 -6
rect 511 -1 513 3
rect 521 -1 523 3
rect 495 -10 497 -6
rect 561 14 563 25
rect 571 23 573 36
rect 656 43 658 48
rect 608 36 610 39
rect 601 34 610 36
rect 618 35 620 39
rect 628 36 630 39
rect 592 26 594 34
rect 601 32 603 34
rect 605 32 610 34
rect 601 30 610 32
rect 626 34 630 36
rect 626 31 628 34
rect 608 26 610 30
rect 622 29 628 31
rect 635 30 637 39
rect 666 40 668 45
rect 676 40 678 45
rect 696 45 698 49
rect 709 47 711 52
rect 716 47 718 52
rect 740 56 765 58
rect 740 48 742 56
rect 753 48 755 52
rect 763 48 765 56
rect 773 51 775 56
rect 780 51 782 56
rect 737 46 742 48
rect 737 43 739 46
rect 656 31 658 34
rect 666 31 668 34
rect 622 27 624 29
rect 626 27 628 29
rect 589 24 602 26
rect 608 24 618 26
rect 622 25 628 27
rect 589 23 591 24
rect 571 21 577 23
rect 571 19 573 21
rect 575 19 577 21
rect 571 17 577 19
rect 585 21 591 23
rect 600 21 602 24
rect 616 21 618 24
rect 626 21 628 25
rect 632 28 638 30
rect 632 26 634 28
rect 636 26 638 28
rect 632 24 638 26
rect 636 21 638 24
rect 656 29 662 31
rect 656 27 658 29
rect 660 27 662 29
rect 656 25 662 27
rect 666 29 672 31
rect 666 27 668 29
rect 670 27 672 29
rect 666 25 672 27
rect 656 22 658 25
rect 585 19 587 21
rect 589 19 591 21
rect 585 17 591 19
rect 571 14 573 17
rect 551 -1 553 3
rect 561 -4 563 1
rect 571 -4 573 1
rect 531 -10 533 -6
rect 616 -1 618 3
rect 626 -1 628 3
rect 600 -10 602 -6
rect 669 15 671 25
rect 676 24 678 34
rect 696 31 698 36
rect 709 31 711 36
rect 696 29 702 31
rect 696 27 698 29
rect 700 27 702 29
rect 696 25 702 27
rect 706 29 712 31
rect 706 27 708 29
rect 710 27 712 29
rect 706 25 712 27
rect 676 22 682 24
rect 676 20 678 22
rect 680 20 682 22
rect 696 21 698 25
rect 676 18 682 20
rect 676 15 678 18
rect 656 -1 658 4
rect 636 -10 638 -6
rect 706 14 708 25
rect 716 23 718 36
rect 801 45 803 49
rect 814 47 816 52
rect 821 47 823 52
rect 845 56 870 58
rect 845 48 847 56
rect 858 48 860 52
rect 868 48 870 56
rect 878 51 880 56
rect 885 51 887 56
rect 753 36 755 39
rect 746 34 755 36
rect 763 35 765 39
rect 773 36 775 39
rect 737 26 739 34
rect 746 32 748 34
rect 750 32 755 34
rect 746 30 755 32
rect 771 34 775 36
rect 771 31 773 34
rect 753 26 755 30
rect 767 29 773 31
rect 780 30 782 39
rect 842 46 847 48
rect 842 43 844 46
rect 801 31 803 36
rect 814 31 816 36
rect 767 27 769 29
rect 771 27 773 29
rect 734 24 747 26
rect 753 24 763 26
rect 767 25 773 27
rect 734 23 736 24
rect 716 21 722 23
rect 716 19 718 21
rect 720 19 722 21
rect 716 17 722 19
rect 730 21 736 23
rect 745 21 747 24
rect 761 21 763 24
rect 771 21 773 25
rect 777 28 783 30
rect 777 26 779 28
rect 781 26 783 28
rect 777 24 783 26
rect 781 21 783 24
rect 801 29 807 31
rect 801 27 803 29
rect 805 27 807 29
rect 801 25 807 27
rect 811 29 817 31
rect 811 27 813 29
rect 815 27 817 29
rect 811 25 817 27
rect 801 21 803 25
rect 730 19 732 21
rect 734 19 736 21
rect 730 17 736 19
rect 716 14 718 17
rect 696 -1 698 3
rect 706 -4 708 1
rect 716 -4 718 1
rect 669 -10 671 -6
rect 676 -10 678 -6
rect 761 -1 763 3
rect 771 -1 773 3
rect 745 -10 747 -6
rect 811 14 813 25
rect 821 23 823 36
rect 906 43 908 48
rect 858 36 860 39
rect 851 34 860 36
rect 868 35 870 39
rect 878 36 880 39
rect 842 26 844 34
rect 851 32 853 34
rect 855 32 860 34
rect 851 30 860 32
rect 876 34 880 36
rect 876 31 878 34
rect 858 26 860 30
rect 872 29 878 31
rect 885 30 887 39
rect 916 40 918 45
rect 926 40 928 45
rect 946 45 948 49
rect 959 47 961 52
rect 966 47 968 52
rect 990 56 1015 58
rect 990 48 992 56
rect 1003 48 1005 52
rect 1013 48 1015 56
rect 1023 51 1025 56
rect 1030 51 1032 56
rect 987 46 992 48
rect 987 43 989 46
rect 906 31 908 34
rect 916 31 918 34
rect 872 27 874 29
rect 876 27 878 29
rect 839 24 852 26
rect 858 24 868 26
rect 872 25 878 27
rect 839 23 841 24
rect 821 21 827 23
rect 821 19 823 21
rect 825 19 827 21
rect 821 17 827 19
rect 835 21 841 23
rect 850 21 852 24
rect 866 21 868 24
rect 876 21 878 25
rect 882 28 888 30
rect 882 26 884 28
rect 886 26 888 28
rect 882 24 888 26
rect 886 21 888 24
rect 906 29 912 31
rect 906 27 908 29
rect 910 27 912 29
rect 906 25 912 27
rect 916 29 922 31
rect 916 27 918 29
rect 920 27 922 29
rect 916 25 922 27
rect 906 22 908 25
rect 835 19 837 21
rect 839 19 841 21
rect 835 17 841 19
rect 821 14 823 17
rect 801 -1 803 3
rect 811 -4 813 1
rect 821 -4 823 1
rect 781 -10 783 -6
rect 866 -1 868 3
rect 876 -1 878 3
rect 850 -10 852 -6
rect 919 15 921 25
rect 926 24 928 34
rect 946 31 948 36
rect 959 31 961 36
rect 946 29 952 31
rect 946 27 948 29
rect 950 27 952 29
rect 946 25 952 27
rect 956 29 962 31
rect 956 27 958 29
rect 960 27 962 29
rect 956 25 962 27
rect 926 22 932 24
rect 926 20 928 22
rect 930 20 932 22
rect 946 21 948 25
rect 926 18 932 20
rect 926 15 928 18
rect 906 -1 908 4
rect 886 -10 888 -6
rect 956 14 958 25
rect 966 23 968 36
rect 1051 45 1053 49
rect 1064 47 1066 52
rect 1071 47 1073 52
rect 1095 56 1120 58
rect 1095 48 1097 56
rect 1108 48 1110 52
rect 1118 48 1120 56
rect 1128 51 1130 56
rect 1135 51 1137 56
rect 1003 36 1005 39
rect 996 34 1005 36
rect 1013 35 1015 39
rect 1023 36 1025 39
rect 987 26 989 34
rect 996 32 998 34
rect 1000 32 1005 34
rect 996 30 1005 32
rect 1021 34 1025 36
rect 1021 31 1023 34
rect 1003 26 1005 30
rect 1017 29 1023 31
rect 1030 30 1032 39
rect 1092 46 1097 48
rect 1092 43 1094 46
rect 1051 31 1053 36
rect 1064 31 1066 36
rect 1017 27 1019 29
rect 1021 27 1023 29
rect 984 24 997 26
rect 1003 24 1013 26
rect 1017 25 1023 27
rect 984 23 986 24
rect 966 21 972 23
rect 966 19 968 21
rect 970 19 972 21
rect 966 17 972 19
rect 980 21 986 23
rect 995 21 997 24
rect 1011 21 1013 24
rect 1021 21 1023 25
rect 1027 28 1033 30
rect 1027 26 1029 28
rect 1031 26 1033 28
rect 1027 24 1033 26
rect 1031 21 1033 24
rect 1051 29 1057 31
rect 1051 27 1053 29
rect 1055 27 1057 29
rect 1051 25 1057 27
rect 1061 29 1067 31
rect 1061 27 1063 29
rect 1065 27 1067 29
rect 1061 25 1067 27
rect 1051 21 1053 25
rect 980 19 982 21
rect 984 19 986 21
rect 980 17 986 19
rect 966 14 968 17
rect 946 -1 948 3
rect 956 -4 958 1
rect 966 -4 968 1
rect 919 -10 921 -6
rect 926 -10 928 -6
rect 1011 -1 1013 3
rect 1021 -1 1023 3
rect 995 -10 997 -6
rect 1061 14 1063 25
rect 1071 23 1073 36
rect 1108 36 1110 39
rect 1101 34 1110 36
rect 1118 35 1120 39
rect 1128 36 1130 39
rect 1092 26 1094 34
rect 1101 32 1103 34
rect 1105 32 1110 34
rect 1101 30 1110 32
rect 1126 34 1130 36
rect 1126 31 1128 34
rect 1108 26 1110 30
rect 1122 29 1128 31
rect 1135 30 1137 39
rect 1122 27 1124 29
rect 1126 27 1128 29
rect 1089 24 1102 26
rect 1108 24 1118 26
rect 1122 25 1128 27
rect 1089 23 1091 24
rect 1071 21 1077 23
rect 1071 19 1073 21
rect 1075 19 1077 21
rect 1071 17 1077 19
rect 1085 21 1091 23
rect 1100 21 1102 24
rect 1116 21 1118 24
rect 1126 21 1128 25
rect 1132 28 1138 30
rect 1132 26 1134 28
rect 1136 26 1138 28
rect 1132 24 1138 26
rect 1136 21 1138 24
rect 1085 19 1087 21
rect 1089 19 1091 21
rect 1085 17 1091 19
rect 1071 14 1073 17
rect 1051 -1 1053 3
rect 1061 -4 1063 1
rect 1071 -4 1073 1
rect 1031 -10 1033 -6
rect 1116 -1 1118 3
rect 1126 -1 1128 3
rect 1100 -10 1102 -6
rect 1136 -10 1138 -6
<< ndif >>
rect 219 343 226 345
rect 219 341 222 343
rect 224 341 226 343
rect 219 335 226 341
rect 259 343 266 345
rect 259 341 262 343
rect 264 341 266 343
rect 201 333 208 335
rect 201 331 203 333
rect 205 331 208 333
rect 201 329 208 331
rect 203 324 208 329
rect 210 324 215 335
rect 217 333 226 335
rect 259 335 266 341
rect 288 343 294 345
rect 288 341 290 343
rect 292 341 294 343
rect 288 339 294 341
rect 241 333 248 335
rect 217 324 228 333
rect 230 331 237 333
rect 230 329 233 331
rect 235 329 237 331
rect 241 331 243 333
rect 245 331 248 333
rect 241 329 248 331
rect 230 327 237 329
rect 230 324 235 327
rect 243 324 248 329
rect 250 324 255 335
rect 257 333 266 335
rect 257 324 268 333
rect 270 331 277 333
rect 270 329 273 331
rect 275 329 277 331
rect 270 327 277 329
rect 288 327 296 339
rect 298 327 303 339
rect 305 336 310 339
rect 371 343 378 345
rect 371 341 374 343
rect 376 341 378 343
rect 305 333 313 336
rect 305 331 308 333
rect 310 331 313 333
rect 305 327 313 331
rect 315 331 323 336
rect 315 329 318 331
rect 320 329 323 331
rect 315 327 323 329
rect 325 334 334 336
rect 371 335 378 341
rect 435 343 442 345
rect 435 341 438 343
rect 440 341 442 343
rect 325 332 330 334
rect 332 332 334 334
rect 325 331 334 332
rect 353 333 360 335
rect 353 331 355 333
rect 357 331 360 333
rect 325 327 339 331
rect 270 324 275 327
rect 334 322 339 327
rect 341 328 346 331
rect 353 329 360 331
rect 341 326 348 328
rect 341 324 344 326
rect 346 324 348 326
rect 355 324 360 329
rect 362 324 367 335
rect 369 333 378 335
rect 435 335 442 341
rect 475 343 482 345
rect 475 341 478 343
rect 480 341 482 343
rect 417 333 424 335
rect 369 324 380 333
rect 382 331 389 333
rect 382 329 385 331
rect 387 329 389 331
rect 417 331 419 333
rect 421 331 424 333
rect 417 329 424 331
rect 382 327 389 329
rect 382 324 387 327
rect 419 324 424 329
rect 426 324 431 335
rect 433 333 442 335
rect 475 335 482 341
rect 504 343 510 345
rect 504 341 506 343
rect 508 341 510 343
rect 504 339 510 341
rect 457 333 464 335
rect 433 324 444 333
rect 446 331 453 333
rect 446 329 449 331
rect 451 329 453 331
rect 457 331 459 333
rect 461 331 464 333
rect 457 329 464 331
rect 446 327 453 329
rect 446 324 451 327
rect 459 324 464 329
rect 466 324 471 335
rect 473 333 482 335
rect 473 324 484 333
rect 486 331 493 333
rect 486 329 489 331
rect 491 329 493 331
rect 486 327 493 329
rect 504 327 512 339
rect 514 327 519 339
rect 521 336 526 339
rect 587 343 594 345
rect 587 341 590 343
rect 592 341 594 343
rect 521 333 529 336
rect 521 331 524 333
rect 526 331 529 333
rect 521 327 529 331
rect 531 331 539 336
rect 531 329 534 331
rect 536 329 539 331
rect 531 327 539 329
rect 541 334 550 336
rect 587 335 594 341
rect 640 343 647 345
rect 640 341 643 343
rect 645 341 647 343
rect 541 332 546 334
rect 548 332 550 334
rect 541 331 550 332
rect 569 333 576 335
rect 569 331 571 333
rect 573 331 576 333
rect 541 327 555 331
rect 486 324 491 327
rect 341 322 348 324
rect 550 322 555 327
rect 557 328 562 331
rect 569 329 576 331
rect 557 326 564 328
rect 557 324 560 326
rect 562 324 564 326
rect 571 324 576 329
rect 578 324 583 335
rect 585 333 594 335
rect 640 335 647 341
rect 680 343 687 345
rect 680 341 683 343
rect 685 341 687 343
rect 622 333 629 335
rect 585 324 596 333
rect 598 331 605 333
rect 598 329 601 331
rect 603 329 605 331
rect 622 331 624 333
rect 626 331 629 333
rect 622 329 629 331
rect 598 327 605 329
rect 598 324 603 327
rect 624 324 629 329
rect 631 324 636 335
rect 638 333 647 335
rect 680 335 687 341
rect 709 343 715 345
rect 709 341 711 343
rect 713 341 715 343
rect 709 339 715 341
rect 662 333 669 335
rect 638 324 649 333
rect 651 331 658 333
rect 651 329 654 331
rect 656 329 658 331
rect 662 331 664 333
rect 666 331 669 333
rect 662 329 669 331
rect 651 327 658 329
rect 651 324 656 327
rect 664 324 669 329
rect 671 324 676 335
rect 678 333 687 335
rect 678 324 689 333
rect 691 331 698 333
rect 691 329 694 331
rect 696 329 698 331
rect 691 327 698 329
rect 709 327 717 339
rect 719 327 724 339
rect 726 336 731 339
rect 792 343 799 345
rect 792 341 795 343
rect 797 341 799 343
rect 726 333 734 336
rect 726 331 729 333
rect 731 331 734 333
rect 726 327 734 331
rect 736 331 744 336
rect 736 329 739 331
rect 741 329 744 331
rect 736 327 744 329
rect 746 334 755 336
rect 792 335 799 341
rect 859 343 866 345
rect 859 341 862 343
rect 864 341 866 343
rect 746 332 751 334
rect 753 332 755 334
rect 746 331 755 332
rect 774 333 781 335
rect 774 331 776 333
rect 778 331 781 333
rect 746 327 760 331
rect 691 324 696 327
rect 557 322 564 324
rect 755 322 760 327
rect 762 328 767 331
rect 774 329 781 331
rect 762 326 769 328
rect 762 324 765 326
rect 767 324 769 326
rect 776 324 781 329
rect 783 324 788 335
rect 790 333 799 335
rect 859 335 866 341
rect 899 343 906 345
rect 899 341 902 343
rect 904 341 906 343
rect 841 333 848 335
rect 790 324 801 333
rect 803 331 810 333
rect 803 329 806 331
rect 808 329 810 331
rect 841 331 843 333
rect 845 331 848 333
rect 841 329 848 331
rect 803 327 810 329
rect 803 324 808 327
rect 843 324 848 329
rect 850 324 855 335
rect 857 333 866 335
rect 899 335 906 341
rect 928 343 934 345
rect 928 341 930 343
rect 932 341 934 343
rect 928 339 934 341
rect 881 333 888 335
rect 857 324 868 333
rect 870 331 877 333
rect 870 329 873 331
rect 875 329 877 331
rect 881 331 883 333
rect 885 331 888 333
rect 881 329 888 331
rect 870 327 877 329
rect 870 324 875 327
rect 883 324 888 329
rect 890 324 895 335
rect 897 333 906 335
rect 897 324 908 333
rect 910 331 917 333
rect 910 329 913 331
rect 915 329 917 331
rect 910 327 917 329
rect 928 327 936 339
rect 938 327 943 339
rect 945 336 950 339
rect 1011 343 1018 345
rect 1011 341 1014 343
rect 1016 341 1018 343
rect 945 333 953 336
rect 945 331 948 333
rect 950 331 953 333
rect 945 327 953 331
rect 955 331 963 336
rect 955 329 958 331
rect 960 329 963 331
rect 955 327 963 329
rect 965 334 974 336
rect 1011 335 1018 341
rect 965 332 970 334
rect 972 332 974 334
rect 965 331 974 332
rect 993 333 1000 335
rect 993 331 995 333
rect 997 331 1000 333
rect 965 327 979 331
rect 910 324 915 327
rect 762 322 769 324
rect 974 322 979 327
rect 981 328 986 331
rect 993 329 1000 331
rect 981 326 988 328
rect 981 324 984 326
rect 986 324 988 326
rect 995 324 1000 329
rect 1002 324 1007 335
rect 1009 333 1018 335
rect 1009 324 1020 333
rect 1022 331 1029 333
rect 1022 329 1025 331
rect 1027 329 1029 331
rect 1022 327 1029 329
rect 1022 324 1027 327
rect 981 322 988 324
rect 322 228 329 230
rect 203 225 208 228
rect 201 223 208 225
rect 201 221 203 223
rect 205 221 208 223
rect 201 219 208 221
rect 210 219 221 228
rect 212 217 221 219
rect 223 217 228 228
rect 230 223 235 228
rect 243 223 248 228
rect 230 221 237 223
rect 230 219 233 221
rect 235 219 237 221
rect 230 217 237 219
rect 241 221 248 223
rect 241 219 243 221
rect 245 219 248 221
rect 241 217 248 219
rect 250 217 255 228
rect 257 219 268 228
rect 270 225 275 228
rect 283 225 288 228
rect 270 223 277 225
rect 270 221 273 223
rect 275 221 277 223
rect 270 219 277 221
rect 281 223 288 225
rect 281 221 283 223
rect 285 221 288 223
rect 281 219 288 221
rect 290 219 301 228
rect 257 217 266 219
rect 212 211 219 217
rect 212 209 214 211
rect 216 209 219 211
rect 212 207 219 209
rect 259 211 266 217
rect 292 217 301 219
rect 303 217 308 228
rect 310 223 315 228
rect 322 226 324 228
rect 326 226 329 228
rect 322 224 329 226
rect 310 221 317 223
rect 324 221 329 224
rect 331 225 336 230
rect 538 228 545 230
rect 419 225 424 228
rect 331 221 345 225
rect 310 219 313 221
rect 315 219 317 221
rect 310 217 317 219
rect 336 220 345 221
rect 336 218 338 220
rect 340 218 345 220
rect 259 209 262 211
rect 264 209 266 211
rect 259 207 266 209
rect 292 211 299 217
rect 336 216 345 218
rect 347 223 355 225
rect 347 221 350 223
rect 352 221 355 223
rect 347 216 355 221
rect 357 221 365 225
rect 357 219 360 221
rect 362 219 365 221
rect 357 216 365 219
rect 292 209 294 211
rect 296 209 299 211
rect 292 207 299 209
rect 360 213 365 216
rect 367 213 372 225
rect 374 213 382 225
rect 417 223 424 225
rect 417 221 419 223
rect 421 221 424 223
rect 417 219 424 221
rect 426 219 437 228
rect 428 217 437 219
rect 439 217 444 228
rect 446 223 451 228
rect 459 223 464 228
rect 446 221 453 223
rect 446 219 449 221
rect 451 219 453 221
rect 446 217 453 219
rect 457 221 464 223
rect 457 219 459 221
rect 461 219 464 221
rect 457 217 464 219
rect 466 217 471 228
rect 473 219 484 228
rect 486 225 491 228
rect 499 225 504 228
rect 486 223 493 225
rect 486 221 489 223
rect 491 221 493 223
rect 486 219 493 221
rect 497 223 504 225
rect 497 221 499 223
rect 501 221 504 223
rect 497 219 504 221
rect 506 219 517 228
rect 473 217 482 219
rect 376 211 382 213
rect 376 209 378 211
rect 380 209 382 211
rect 376 207 382 209
rect 428 211 435 217
rect 428 209 430 211
rect 432 209 435 211
rect 428 207 435 209
rect 475 211 482 217
rect 508 217 517 219
rect 519 217 524 228
rect 526 223 531 228
rect 538 226 540 228
rect 542 226 545 228
rect 538 224 545 226
rect 526 221 533 223
rect 540 221 545 224
rect 547 225 552 230
rect 743 228 750 230
rect 624 225 629 228
rect 547 221 561 225
rect 526 219 529 221
rect 531 219 533 221
rect 526 217 533 219
rect 552 220 561 221
rect 552 218 554 220
rect 556 218 561 220
rect 475 209 478 211
rect 480 209 482 211
rect 475 207 482 209
rect 508 211 515 217
rect 552 216 561 218
rect 563 223 571 225
rect 563 221 566 223
rect 568 221 571 223
rect 563 216 571 221
rect 573 221 581 225
rect 573 219 576 221
rect 578 219 581 221
rect 573 216 581 219
rect 508 209 510 211
rect 512 209 515 211
rect 508 207 515 209
rect 576 213 581 216
rect 583 213 588 225
rect 590 213 598 225
rect 622 223 629 225
rect 622 221 624 223
rect 626 221 629 223
rect 622 219 629 221
rect 631 219 642 228
rect 633 217 642 219
rect 644 217 649 228
rect 651 223 656 228
rect 664 223 669 228
rect 651 221 658 223
rect 651 219 654 221
rect 656 219 658 221
rect 651 217 658 219
rect 662 221 669 223
rect 662 219 664 221
rect 666 219 669 221
rect 662 217 669 219
rect 671 217 676 228
rect 678 219 689 228
rect 691 225 696 228
rect 704 225 709 228
rect 691 223 698 225
rect 691 221 694 223
rect 696 221 698 223
rect 691 219 698 221
rect 702 223 709 225
rect 702 221 704 223
rect 706 221 709 223
rect 702 219 709 221
rect 711 219 722 228
rect 678 217 687 219
rect 592 211 598 213
rect 592 209 594 211
rect 596 209 598 211
rect 592 207 598 209
rect 633 211 640 217
rect 633 209 635 211
rect 637 209 640 211
rect 633 207 640 209
rect 680 211 687 217
rect 713 217 722 219
rect 724 217 729 228
rect 731 223 736 228
rect 743 226 745 228
rect 747 226 750 228
rect 743 224 750 226
rect 731 221 738 223
rect 745 221 750 224
rect 752 225 757 230
rect 962 228 969 230
rect 843 225 848 228
rect 752 221 766 225
rect 731 219 734 221
rect 736 219 738 221
rect 731 217 738 219
rect 757 220 766 221
rect 757 218 759 220
rect 761 218 766 220
rect 680 209 683 211
rect 685 209 687 211
rect 680 207 687 209
rect 713 211 720 217
rect 757 216 766 218
rect 768 223 776 225
rect 768 221 771 223
rect 773 221 776 223
rect 768 216 776 221
rect 778 221 786 225
rect 778 219 781 221
rect 783 219 786 221
rect 778 216 786 219
rect 713 209 715 211
rect 717 209 720 211
rect 713 207 720 209
rect 781 213 786 216
rect 788 213 793 225
rect 795 213 803 225
rect 841 223 848 225
rect 841 221 843 223
rect 845 221 848 223
rect 841 219 848 221
rect 850 219 861 228
rect 852 217 861 219
rect 863 217 868 228
rect 870 223 875 228
rect 883 223 888 228
rect 870 221 877 223
rect 870 219 873 221
rect 875 219 877 221
rect 870 217 877 219
rect 881 221 888 223
rect 881 219 883 221
rect 885 219 888 221
rect 881 217 888 219
rect 890 217 895 228
rect 897 219 908 228
rect 910 225 915 228
rect 923 225 928 228
rect 910 223 917 225
rect 910 221 913 223
rect 915 221 917 223
rect 910 219 917 221
rect 921 223 928 225
rect 921 221 923 223
rect 925 221 928 223
rect 921 219 928 221
rect 930 219 941 228
rect 897 217 906 219
rect 797 211 803 213
rect 797 209 799 211
rect 801 209 803 211
rect 797 207 803 209
rect 852 211 859 217
rect 852 209 854 211
rect 856 209 859 211
rect 852 207 859 209
rect 899 211 906 217
rect 932 217 941 219
rect 943 217 948 228
rect 950 223 955 228
rect 962 226 964 228
rect 966 226 969 228
rect 962 224 969 226
rect 950 221 957 223
rect 964 221 969 224
rect 971 225 976 230
rect 1086 228 1093 230
rect 1047 225 1052 228
rect 971 221 985 225
rect 950 219 953 221
rect 955 219 957 221
rect 950 217 957 219
rect 976 220 985 221
rect 976 218 978 220
rect 980 218 985 220
rect 899 209 902 211
rect 904 209 906 211
rect 899 207 906 209
rect 932 211 939 217
rect 976 216 985 218
rect 987 223 995 225
rect 987 221 990 223
rect 992 221 995 223
rect 987 216 995 221
rect 997 221 1005 225
rect 997 219 1000 221
rect 1002 219 1005 221
rect 997 216 1005 219
rect 932 209 934 211
rect 936 209 939 211
rect 932 207 939 209
rect 1000 213 1005 216
rect 1007 213 1012 225
rect 1014 213 1022 225
rect 1045 223 1052 225
rect 1045 221 1047 223
rect 1049 221 1052 223
rect 1045 219 1052 221
rect 1054 219 1065 228
rect 1056 217 1065 219
rect 1067 217 1072 228
rect 1074 223 1079 228
rect 1086 226 1088 228
rect 1090 226 1093 228
rect 1086 224 1093 226
rect 1074 221 1081 223
rect 1088 221 1093 224
rect 1095 225 1100 230
rect 1095 221 1109 225
rect 1074 219 1077 221
rect 1079 219 1081 221
rect 1074 217 1081 219
rect 1100 220 1109 221
rect 1100 218 1102 220
rect 1104 218 1109 220
rect 1016 211 1022 213
rect 1016 209 1018 211
rect 1020 209 1022 211
rect 1016 207 1022 209
rect 1056 211 1063 217
rect 1100 216 1109 218
rect 1111 223 1119 225
rect 1111 221 1114 223
rect 1116 221 1119 223
rect 1111 216 1119 221
rect 1121 221 1129 225
rect 1121 219 1124 221
rect 1126 219 1129 221
rect 1121 216 1129 219
rect 1056 209 1058 211
rect 1060 209 1063 211
rect 1056 207 1063 209
rect 1124 213 1129 216
rect 1131 213 1136 225
rect 1138 213 1146 225
rect 1140 211 1146 213
rect 1140 209 1142 211
rect 1144 209 1146 211
rect 1140 207 1146 209
rect 162 195 168 197
rect 162 193 164 195
rect 166 193 168 195
rect 162 191 168 193
rect 181 195 187 197
rect 202 199 209 201
rect 202 197 204 199
rect 206 197 209 199
rect 181 193 183 195
rect 185 193 187 195
rect 181 191 187 193
rect 162 187 166 191
rect 153 184 158 187
rect 151 182 158 184
rect 151 180 153 182
rect 155 180 158 182
rect 151 178 158 180
rect 160 184 166 187
rect 182 184 187 191
rect 202 191 209 197
rect 286 199 292 201
rect 286 197 288 199
rect 290 197 292 199
rect 286 195 292 197
rect 307 199 314 201
rect 307 197 309 199
rect 311 197 314 199
rect 270 192 275 195
rect 202 189 211 191
rect 160 178 168 184
rect 170 182 178 184
rect 170 180 173 182
rect 175 180 178 182
rect 170 178 178 180
rect 180 178 187 184
rect 191 187 198 189
rect 191 185 193 187
rect 195 185 198 187
rect 191 183 198 185
rect 193 180 198 183
rect 200 180 211 189
rect 213 180 218 191
rect 220 189 227 191
rect 220 187 223 189
rect 225 187 227 189
rect 246 190 255 192
rect 246 188 248 190
rect 250 188 255 190
rect 246 187 255 188
rect 220 185 227 187
rect 220 180 225 185
rect 234 184 239 187
rect 232 182 239 184
rect 232 180 234 182
rect 236 180 239 182
rect 232 178 239 180
rect 241 183 255 187
rect 257 187 265 192
rect 257 185 260 187
rect 262 185 265 187
rect 257 183 265 185
rect 267 189 275 192
rect 267 187 270 189
rect 272 187 275 189
rect 267 183 275 187
rect 277 183 282 195
rect 284 183 292 195
rect 307 191 314 197
rect 391 199 397 201
rect 391 197 393 199
rect 395 197 397 199
rect 391 195 397 197
rect 412 195 418 197
rect 375 192 380 195
rect 307 189 316 191
rect 296 187 303 189
rect 296 185 298 187
rect 300 185 303 187
rect 296 183 303 185
rect 241 178 246 183
rect 298 180 303 183
rect 305 180 316 189
rect 318 180 323 191
rect 325 189 332 191
rect 325 187 328 189
rect 330 187 332 189
rect 351 190 360 192
rect 351 188 353 190
rect 355 188 360 190
rect 351 187 360 188
rect 325 185 332 187
rect 325 180 330 185
rect 339 184 344 187
rect 337 182 344 184
rect 337 180 339 182
rect 341 180 344 182
rect 337 178 344 180
rect 346 183 360 187
rect 362 187 370 192
rect 362 185 365 187
rect 367 185 370 187
rect 362 183 370 185
rect 372 189 380 192
rect 372 187 375 189
rect 377 187 380 189
rect 372 183 380 187
rect 382 183 387 195
rect 389 183 397 195
rect 412 193 414 195
rect 416 193 418 195
rect 412 191 418 193
rect 431 195 437 197
rect 452 199 459 201
rect 452 197 454 199
rect 456 197 459 199
rect 431 193 433 195
rect 435 193 437 195
rect 431 191 437 193
rect 412 187 416 191
rect 403 184 408 187
rect 346 178 351 183
rect 401 182 408 184
rect 401 180 403 182
rect 405 180 408 182
rect 401 178 408 180
rect 410 184 416 187
rect 432 184 437 191
rect 452 191 459 197
rect 536 199 542 201
rect 536 197 538 199
rect 540 197 542 199
rect 536 195 542 197
rect 557 199 564 201
rect 557 197 559 199
rect 561 197 564 199
rect 520 192 525 195
rect 452 189 461 191
rect 410 178 418 184
rect 420 182 428 184
rect 420 180 423 182
rect 425 180 428 182
rect 420 178 428 180
rect 430 178 437 184
rect 441 187 448 189
rect 441 185 443 187
rect 445 185 448 187
rect 441 183 448 185
rect 443 180 448 183
rect 450 180 461 189
rect 463 180 468 191
rect 470 189 477 191
rect 470 187 473 189
rect 475 187 477 189
rect 496 190 505 192
rect 496 188 498 190
rect 500 188 505 190
rect 496 187 505 188
rect 470 185 477 187
rect 470 180 475 185
rect 484 184 489 187
rect 482 182 489 184
rect 482 180 484 182
rect 486 180 489 182
rect 482 178 489 180
rect 491 183 505 187
rect 507 187 515 192
rect 507 185 510 187
rect 512 185 515 187
rect 507 183 515 185
rect 517 189 525 192
rect 517 187 520 189
rect 522 187 525 189
rect 517 183 525 187
rect 527 183 532 195
rect 534 183 542 195
rect 557 191 564 197
rect 641 199 647 201
rect 641 197 643 199
rect 645 197 647 199
rect 641 195 647 197
rect 662 195 668 197
rect 625 192 630 195
rect 557 189 566 191
rect 546 187 553 189
rect 546 185 548 187
rect 550 185 553 187
rect 546 183 553 185
rect 491 178 496 183
rect 548 180 553 183
rect 555 180 566 189
rect 568 180 573 191
rect 575 189 582 191
rect 575 187 578 189
rect 580 187 582 189
rect 601 190 610 192
rect 601 188 603 190
rect 605 188 610 190
rect 601 187 610 188
rect 575 185 582 187
rect 575 180 580 185
rect 589 184 594 187
rect 587 182 594 184
rect 587 180 589 182
rect 591 180 594 182
rect 587 178 594 180
rect 596 183 610 187
rect 612 187 620 192
rect 612 185 615 187
rect 617 185 620 187
rect 612 183 620 185
rect 622 189 630 192
rect 622 187 625 189
rect 627 187 630 189
rect 622 183 630 187
rect 632 183 637 195
rect 639 183 647 195
rect 662 193 664 195
rect 666 193 668 195
rect 662 191 668 193
rect 681 195 687 197
rect 702 199 709 201
rect 702 197 704 199
rect 706 197 709 199
rect 681 193 683 195
rect 685 193 687 195
rect 681 191 687 193
rect 662 187 666 191
rect 653 184 658 187
rect 596 178 601 183
rect 651 182 658 184
rect 651 180 653 182
rect 655 180 658 182
rect 651 178 658 180
rect 660 184 666 187
rect 682 184 687 191
rect 702 191 709 197
rect 786 199 792 201
rect 786 197 788 199
rect 790 197 792 199
rect 786 195 792 197
rect 807 199 814 201
rect 807 197 809 199
rect 811 197 814 199
rect 770 192 775 195
rect 702 189 711 191
rect 660 178 668 184
rect 670 182 678 184
rect 670 180 673 182
rect 675 180 678 182
rect 670 178 678 180
rect 680 178 687 184
rect 691 187 698 189
rect 691 185 693 187
rect 695 185 698 187
rect 691 183 698 185
rect 693 180 698 183
rect 700 180 711 189
rect 713 180 718 191
rect 720 189 727 191
rect 720 187 723 189
rect 725 187 727 189
rect 746 190 755 192
rect 746 188 748 190
rect 750 188 755 190
rect 746 187 755 188
rect 720 185 727 187
rect 720 180 725 185
rect 734 184 739 187
rect 732 182 739 184
rect 732 180 734 182
rect 736 180 739 182
rect 732 178 739 180
rect 741 183 755 187
rect 757 187 765 192
rect 757 185 760 187
rect 762 185 765 187
rect 757 183 765 185
rect 767 189 775 192
rect 767 187 770 189
rect 772 187 775 189
rect 767 183 775 187
rect 777 183 782 195
rect 784 183 792 195
rect 807 191 814 197
rect 891 199 897 201
rect 891 197 893 199
rect 895 197 897 199
rect 891 195 897 197
rect 912 195 918 197
rect 875 192 880 195
rect 807 189 816 191
rect 796 187 803 189
rect 796 185 798 187
rect 800 185 803 187
rect 796 183 803 185
rect 741 178 746 183
rect 798 180 803 183
rect 805 180 816 189
rect 818 180 823 191
rect 825 189 832 191
rect 825 187 828 189
rect 830 187 832 189
rect 851 190 860 192
rect 851 188 853 190
rect 855 188 860 190
rect 851 187 860 188
rect 825 185 832 187
rect 825 180 830 185
rect 839 184 844 187
rect 837 182 844 184
rect 837 180 839 182
rect 841 180 844 182
rect 837 178 844 180
rect 846 183 860 187
rect 862 187 870 192
rect 862 185 865 187
rect 867 185 870 187
rect 862 183 870 185
rect 872 189 880 192
rect 872 187 875 189
rect 877 187 880 189
rect 872 183 880 187
rect 882 183 887 195
rect 889 183 897 195
rect 912 193 914 195
rect 916 193 918 195
rect 912 191 918 193
rect 931 195 937 197
rect 952 199 959 201
rect 952 197 954 199
rect 956 197 959 199
rect 931 193 933 195
rect 935 193 937 195
rect 931 191 937 193
rect 912 187 916 191
rect 903 184 908 187
rect 846 178 851 183
rect 901 182 908 184
rect 901 180 903 182
rect 905 180 908 182
rect 901 178 908 180
rect 910 184 916 187
rect 932 184 937 191
rect 952 191 959 197
rect 1036 199 1042 201
rect 1036 197 1038 199
rect 1040 197 1042 199
rect 1036 195 1042 197
rect 1057 199 1064 201
rect 1057 197 1059 199
rect 1061 197 1064 199
rect 1020 192 1025 195
rect 952 189 961 191
rect 910 178 918 184
rect 920 182 928 184
rect 920 180 923 182
rect 925 180 928 182
rect 920 178 928 180
rect 930 178 937 184
rect 941 187 948 189
rect 941 185 943 187
rect 945 185 948 187
rect 941 183 948 185
rect 943 180 948 183
rect 950 180 961 189
rect 963 180 968 191
rect 970 189 977 191
rect 970 187 973 189
rect 975 187 977 189
rect 996 190 1005 192
rect 996 188 998 190
rect 1000 188 1005 190
rect 996 187 1005 188
rect 970 185 977 187
rect 970 180 975 185
rect 984 184 989 187
rect 982 182 989 184
rect 982 180 984 182
rect 986 180 989 182
rect 982 178 989 180
rect 991 183 1005 187
rect 1007 187 1015 192
rect 1007 185 1010 187
rect 1012 185 1015 187
rect 1007 183 1015 185
rect 1017 189 1025 192
rect 1017 187 1020 189
rect 1022 187 1025 189
rect 1017 183 1025 187
rect 1027 183 1032 195
rect 1034 183 1042 195
rect 1057 191 1064 197
rect 1141 199 1147 201
rect 1141 197 1143 199
rect 1145 197 1147 199
rect 1141 195 1147 197
rect 1125 192 1130 195
rect 1057 189 1066 191
rect 1046 187 1053 189
rect 1046 185 1048 187
rect 1050 185 1053 187
rect 1046 183 1053 185
rect 991 178 996 183
rect 1048 180 1053 183
rect 1055 180 1066 189
rect 1068 180 1073 191
rect 1075 189 1082 191
rect 1075 187 1078 189
rect 1080 187 1082 189
rect 1101 190 1110 192
rect 1101 188 1103 190
rect 1105 188 1110 190
rect 1101 187 1110 188
rect 1075 185 1082 187
rect 1075 180 1080 185
rect 1089 184 1094 187
rect 1087 182 1094 184
rect 1087 180 1089 182
rect 1091 180 1094 182
rect 1087 178 1094 180
rect 1096 183 1110 187
rect 1112 187 1120 192
rect 1112 185 1115 187
rect 1117 185 1120 187
rect 1112 183 1120 185
rect 1122 189 1130 192
rect 1122 187 1125 189
rect 1127 187 1130 189
rect 1122 183 1130 187
rect 1132 183 1137 195
rect 1139 183 1147 195
rect 1096 178 1101 183
rect 150 84 157 86
rect 150 82 152 84
rect 154 82 157 84
rect 150 80 157 82
rect 152 77 157 80
rect 159 80 167 86
rect 169 84 177 86
rect 169 82 172 84
rect 174 82 177 84
rect 169 80 177 82
rect 179 80 186 86
rect 231 84 238 86
rect 192 81 197 84
rect 159 77 165 80
rect 161 73 165 77
rect 181 73 186 80
rect 190 79 197 81
rect 190 77 192 79
rect 194 77 197 79
rect 190 75 197 77
rect 199 75 210 84
rect 161 71 167 73
rect 161 69 163 71
rect 165 69 167 71
rect 161 67 167 69
rect 180 71 186 73
rect 201 73 210 75
rect 212 73 217 84
rect 219 79 224 84
rect 231 82 233 84
rect 235 82 238 84
rect 231 80 238 82
rect 219 77 226 79
rect 233 77 238 80
rect 240 81 245 86
rect 336 84 343 86
rect 297 81 302 84
rect 240 77 254 81
rect 219 75 222 77
rect 224 75 226 77
rect 219 73 226 75
rect 245 76 254 77
rect 245 74 247 76
rect 249 74 254 76
rect 180 69 182 71
rect 184 69 186 71
rect 180 67 186 69
rect 201 67 208 73
rect 245 72 254 74
rect 256 79 264 81
rect 256 77 259 79
rect 261 77 264 79
rect 256 72 264 77
rect 266 77 274 81
rect 266 75 269 77
rect 271 75 274 77
rect 266 72 274 75
rect 201 65 203 67
rect 205 65 208 67
rect 201 63 208 65
rect 269 69 274 72
rect 276 69 281 81
rect 283 69 291 81
rect 295 79 302 81
rect 295 77 297 79
rect 299 77 302 79
rect 295 75 302 77
rect 304 75 315 84
rect 306 73 315 75
rect 317 73 322 84
rect 324 79 329 84
rect 336 82 338 84
rect 340 82 343 84
rect 336 80 343 82
rect 324 77 331 79
rect 338 77 343 80
rect 345 81 350 86
rect 400 84 407 86
rect 400 82 402 84
rect 404 82 407 84
rect 345 77 359 81
rect 324 75 327 77
rect 329 75 331 77
rect 324 73 331 75
rect 350 76 359 77
rect 350 74 352 76
rect 354 74 359 76
rect 285 67 291 69
rect 285 65 287 67
rect 289 65 291 67
rect 285 63 291 65
rect 306 67 313 73
rect 350 72 359 74
rect 361 79 369 81
rect 361 77 364 79
rect 366 77 369 79
rect 361 72 369 77
rect 371 77 379 81
rect 371 75 374 77
rect 376 75 379 77
rect 371 72 379 75
rect 306 65 308 67
rect 310 65 313 67
rect 306 63 313 65
rect 374 69 379 72
rect 381 69 386 81
rect 388 69 396 81
rect 400 80 407 82
rect 402 77 407 80
rect 409 80 417 86
rect 419 84 427 86
rect 419 82 422 84
rect 424 82 427 84
rect 419 80 427 82
rect 429 80 436 86
rect 481 84 488 86
rect 442 81 447 84
rect 409 77 415 80
rect 411 73 415 77
rect 431 73 436 80
rect 440 79 447 81
rect 440 77 442 79
rect 444 77 447 79
rect 440 75 447 77
rect 449 75 460 84
rect 411 71 417 73
rect 411 69 413 71
rect 415 69 417 71
rect 390 67 396 69
rect 390 65 392 67
rect 394 65 396 67
rect 390 63 396 65
rect 411 67 417 69
rect 430 71 436 73
rect 451 73 460 75
rect 462 73 467 84
rect 469 79 474 84
rect 481 82 483 84
rect 485 82 488 84
rect 481 80 488 82
rect 469 77 476 79
rect 483 77 488 80
rect 490 81 495 86
rect 586 84 593 86
rect 547 81 552 84
rect 490 77 504 81
rect 469 75 472 77
rect 474 75 476 77
rect 469 73 476 75
rect 495 76 504 77
rect 495 74 497 76
rect 499 74 504 76
rect 430 69 432 71
rect 434 69 436 71
rect 430 67 436 69
rect 451 67 458 73
rect 495 72 504 74
rect 506 79 514 81
rect 506 77 509 79
rect 511 77 514 79
rect 506 72 514 77
rect 516 77 524 81
rect 516 75 519 77
rect 521 75 524 77
rect 516 72 524 75
rect 451 65 453 67
rect 455 65 458 67
rect 451 63 458 65
rect 519 69 524 72
rect 526 69 531 81
rect 533 69 541 81
rect 545 79 552 81
rect 545 77 547 79
rect 549 77 552 79
rect 545 75 552 77
rect 554 75 565 84
rect 556 73 565 75
rect 567 73 572 84
rect 574 79 579 84
rect 586 82 588 84
rect 590 82 593 84
rect 586 80 593 82
rect 574 77 581 79
rect 588 77 593 80
rect 595 81 600 86
rect 650 84 657 86
rect 650 82 652 84
rect 654 82 657 84
rect 595 77 609 81
rect 574 75 577 77
rect 579 75 581 77
rect 574 73 581 75
rect 600 76 609 77
rect 600 74 602 76
rect 604 74 609 76
rect 535 67 541 69
rect 535 65 537 67
rect 539 65 541 67
rect 535 63 541 65
rect 556 67 563 73
rect 600 72 609 74
rect 611 79 619 81
rect 611 77 614 79
rect 616 77 619 79
rect 611 72 619 77
rect 621 77 629 81
rect 621 75 624 77
rect 626 75 629 77
rect 621 72 629 75
rect 556 65 558 67
rect 560 65 563 67
rect 556 63 563 65
rect 624 69 629 72
rect 631 69 636 81
rect 638 69 646 81
rect 650 80 657 82
rect 652 77 657 80
rect 659 80 667 86
rect 669 84 677 86
rect 669 82 672 84
rect 674 82 677 84
rect 669 80 677 82
rect 679 80 686 86
rect 731 84 738 86
rect 692 81 697 84
rect 659 77 665 80
rect 661 73 665 77
rect 681 73 686 80
rect 690 79 697 81
rect 690 77 692 79
rect 694 77 697 79
rect 690 75 697 77
rect 699 75 710 84
rect 661 71 667 73
rect 661 69 663 71
rect 665 69 667 71
rect 640 67 646 69
rect 640 65 642 67
rect 644 65 646 67
rect 640 63 646 65
rect 661 67 667 69
rect 680 71 686 73
rect 701 73 710 75
rect 712 73 717 84
rect 719 79 724 84
rect 731 82 733 84
rect 735 82 738 84
rect 731 80 738 82
rect 719 77 726 79
rect 733 77 738 80
rect 740 81 745 86
rect 836 84 843 86
rect 797 81 802 84
rect 740 77 754 81
rect 719 75 722 77
rect 724 75 726 77
rect 719 73 726 75
rect 745 76 754 77
rect 745 74 747 76
rect 749 74 754 76
rect 680 69 682 71
rect 684 69 686 71
rect 680 67 686 69
rect 701 67 708 73
rect 745 72 754 74
rect 756 79 764 81
rect 756 77 759 79
rect 761 77 764 79
rect 756 72 764 77
rect 766 77 774 81
rect 766 75 769 77
rect 771 75 774 77
rect 766 72 774 75
rect 701 65 703 67
rect 705 65 708 67
rect 701 63 708 65
rect 769 69 774 72
rect 776 69 781 81
rect 783 69 791 81
rect 795 79 802 81
rect 795 77 797 79
rect 799 77 802 79
rect 795 75 802 77
rect 804 75 815 84
rect 806 73 815 75
rect 817 73 822 84
rect 824 79 829 84
rect 836 82 838 84
rect 840 82 843 84
rect 836 80 843 82
rect 824 77 831 79
rect 838 77 843 80
rect 845 81 850 86
rect 900 84 907 86
rect 900 82 902 84
rect 904 82 907 84
rect 845 77 859 81
rect 824 75 827 77
rect 829 75 831 77
rect 824 73 831 75
rect 850 76 859 77
rect 850 74 852 76
rect 854 74 859 76
rect 785 67 791 69
rect 785 65 787 67
rect 789 65 791 67
rect 785 63 791 65
rect 806 67 813 73
rect 850 72 859 74
rect 861 79 869 81
rect 861 77 864 79
rect 866 77 869 79
rect 861 72 869 77
rect 871 77 879 81
rect 871 75 874 77
rect 876 75 879 77
rect 871 72 879 75
rect 806 65 808 67
rect 810 65 813 67
rect 806 63 813 65
rect 874 69 879 72
rect 881 69 886 81
rect 888 69 896 81
rect 900 80 907 82
rect 902 77 907 80
rect 909 80 917 86
rect 919 84 927 86
rect 919 82 922 84
rect 924 82 927 84
rect 919 80 927 82
rect 929 80 936 86
rect 981 84 988 86
rect 942 81 947 84
rect 909 77 915 80
rect 911 73 915 77
rect 931 73 936 80
rect 940 79 947 81
rect 940 77 942 79
rect 944 77 947 79
rect 940 75 947 77
rect 949 75 960 84
rect 911 71 917 73
rect 911 69 913 71
rect 915 69 917 71
rect 890 67 896 69
rect 890 65 892 67
rect 894 65 896 67
rect 890 63 896 65
rect 911 67 917 69
rect 930 71 936 73
rect 951 73 960 75
rect 962 73 967 84
rect 969 79 974 84
rect 981 82 983 84
rect 985 82 988 84
rect 981 80 988 82
rect 969 77 976 79
rect 983 77 988 80
rect 990 81 995 86
rect 1086 84 1093 86
rect 1047 81 1052 84
rect 990 77 1004 81
rect 969 75 972 77
rect 974 75 976 77
rect 969 73 976 75
rect 995 76 1004 77
rect 995 74 997 76
rect 999 74 1004 76
rect 930 69 932 71
rect 934 69 936 71
rect 930 67 936 69
rect 951 67 958 73
rect 995 72 1004 74
rect 1006 79 1014 81
rect 1006 77 1009 79
rect 1011 77 1014 79
rect 1006 72 1014 77
rect 1016 77 1024 81
rect 1016 75 1019 77
rect 1021 75 1024 77
rect 1016 72 1024 75
rect 951 65 953 67
rect 955 65 958 67
rect 951 63 958 65
rect 1019 69 1024 72
rect 1026 69 1031 81
rect 1033 69 1041 81
rect 1045 79 1052 81
rect 1045 77 1047 79
rect 1049 77 1052 79
rect 1045 75 1052 77
rect 1054 75 1065 84
rect 1056 73 1065 75
rect 1067 73 1072 84
rect 1074 79 1079 84
rect 1086 82 1088 84
rect 1090 82 1093 84
rect 1086 80 1093 82
rect 1074 77 1081 79
rect 1088 77 1093 80
rect 1095 81 1100 86
rect 1095 77 1109 81
rect 1074 75 1077 77
rect 1079 75 1081 77
rect 1074 73 1081 75
rect 1100 76 1109 77
rect 1100 74 1102 76
rect 1104 74 1109 76
rect 1035 67 1041 69
rect 1035 65 1037 67
rect 1039 65 1041 67
rect 1035 63 1041 65
rect 1056 67 1063 73
rect 1100 72 1109 74
rect 1111 79 1119 81
rect 1111 77 1114 79
rect 1116 77 1119 79
rect 1111 72 1119 77
rect 1121 77 1129 81
rect 1121 75 1124 77
rect 1126 75 1129 77
rect 1121 72 1129 75
rect 1056 65 1058 67
rect 1060 65 1063 67
rect 1056 63 1063 65
rect 1124 69 1129 72
rect 1131 69 1136 81
rect 1138 69 1146 81
rect 1140 67 1146 69
rect 1140 65 1142 67
rect 1144 65 1146 67
rect 1140 63 1146 65
rect 160 51 166 53
rect 160 49 162 51
rect 164 49 166 51
rect 160 47 166 49
rect 179 51 185 53
rect 200 55 207 57
rect 200 53 202 55
rect 204 53 207 55
rect 179 49 181 51
rect 183 49 185 51
rect 179 47 185 49
rect 160 43 164 47
rect 151 40 156 43
rect 149 38 156 40
rect 149 36 151 38
rect 153 36 156 38
rect 149 34 156 36
rect 158 40 164 43
rect 180 40 185 47
rect 200 47 207 53
rect 284 55 290 57
rect 284 53 286 55
rect 288 53 290 55
rect 284 51 290 53
rect 305 55 312 57
rect 305 53 307 55
rect 309 53 312 55
rect 268 48 273 51
rect 200 45 209 47
rect 158 34 166 40
rect 168 38 176 40
rect 168 36 171 38
rect 173 36 176 38
rect 168 34 176 36
rect 178 34 185 40
rect 189 43 196 45
rect 189 41 191 43
rect 193 41 196 43
rect 189 39 196 41
rect 191 36 196 39
rect 198 36 209 45
rect 211 36 216 47
rect 218 45 225 47
rect 218 43 221 45
rect 223 43 225 45
rect 244 46 253 48
rect 244 44 246 46
rect 248 44 253 46
rect 244 43 253 44
rect 218 41 225 43
rect 218 36 223 41
rect 232 40 237 43
rect 230 38 237 40
rect 230 36 232 38
rect 234 36 237 38
rect 230 34 237 36
rect 239 39 253 43
rect 255 43 263 48
rect 255 41 258 43
rect 260 41 263 43
rect 255 39 263 41
rect 265 45 273 48
rect 265 43 268 45
rect 270 43 273 45
rect 265 39 273 43
rect 275 39 280 51
rect 282 39 290 51
rect 305 47 312 53
rect 389 55 395 57
rect 389 53 391 55
rect 393 53 395 55
rect 389 51 395 53
rect 410 51 416 53
rect 373 48 378 51
rect 305 45 314 47
rect 294 43 301 45
rect 294 41 296 43
rect 298 41 301 43
rect 294 39 301 41
rect 239 34 244 39
rect 296 36 301 39
rect 303 36 314 45
rect 316 36 321 47
rect 323 45 330 47
rect 323 43 326 45
rect 328 43 330 45
rect 349 46 358 48
rect 349 44 351 46
rect 353 44 358 46
rect 349 43 358 44
rect 323 41 330 43
rect 323 36 328 41
rect 337 40 342 43
rect 335 38 342 40
rect 335 36 337 38
rect 339 36 342 38
rect 335 34 342 36
rect 344 39 358 43
rect 360 43 368 48
rect 360 41 363 43
rect 365 41 368 43
rect 360 39 368 41
rect 370 45 378 48
rect 370 43 373 45
rect 375 43 378 45
rect 370 39 378 43
rect 380 39 385 51
rect 387 39 395 51
rect 410 49 412 51
rect 414 49 416 51
rect 410 47 416 49
rect 429 51 435 53
rect 450 55 457 57
rect 450 53 452 55
rect 454 53 457 55
rect 429 49 431 51
rect 433 49 435 51
rect 429 47 435 49
rect 410 43 414 47
rect 401 40 406 43
rect 344 34 349 39
rect 399 38 406 40
rect 399 36 401 38
rect 403 36 406 38
rect 399 34 406 36
rect 408 40 414 43
rect 430 40 435 47
rect 450 47 457 53
rect 534 55 540 57
rect 534 53 536 55
rect 538 53 540 55
rect 534 51 540 53
rect 555 55 562 57
rect 555 53 557 55
rect 559 53 562 55
rect 518 48 523 51
rect 450 45 459 47
rect 408 34 416 40
rect 418 38 426 40
rect 418 36 421 38
rect 423 36 426 38
rect 418 34 426 36
rect 428 34 435 40
rect 439 43 446 45
rect 439 41 441 43
rect 443 41 446 43
rect 439 39 446 41
rect 441 36 446 39
rect 448 36 459 45
rect 461 36 466 47
rect 468 45 475 47
rect 468 43 471 45
rect 473 43 475 45
rect 494 46 503 48
rect 494 44 496 46
rect 498 44 503 46
rect 494 43 503 44
rect 468 41 475 43
rect 468 36 473 41
rect 482 40 487 43
rect 480 38 487 40
rect 480 36 482 38
rect 484 36 487 38
rect 480 34 487 36
rect 489 39 503 43
rect 505 43 513 48
rect 505 41 508 43
rect 510 41 513 43
rect 505 39 513 41
rect 515 45 523 48
rect 515 43 518 45
rect 520 43 523 45
rect 515 39 523 43
rect 525 39 530 51
rect 532 39 540 51
rect 555 47 562 53
rect 639 55 645 57
rect 639 53 641 55
rect 643 53 645 55
rect 639 51 645 53
rect 660 51 666 53
rect 623 48 628 51
rect 555 45 564 47
rect 544 43 551 45
rect 544 41 546 43
rect 548 41 551 43
rect 544 39 551 41
rect 489 34 494 39
rect 546 36 551 39
rect 553 36 564 45
rect 566 36 571 47
rect 573 45 580 47
rect 573 43 576 45
rect 578 43 580 45
rect 599 46 608 48
rect 599 44 601 46
rect 603 44 608 46
rect 599 43 608 44
rect 573 41 580 43
rect 573 36 578 41
rect 587 40 592 43
rect 585 38 592 40
rect 585 36 587 38
rect 589 36 592 38
rect 585 34 592 36
rect 594 39 608 43
rect 610 43 618 48
rect 610 41 613 43
rect 615 41 618 43
rect 610 39 618 41
rect 620 45 628 48
rect 620 43 623 45
rect 625 43 628 45
rect 620 39 628 43
rect 630 39 635 51
rect 637 39 645 51
rect 660 49 662 51
rect 664 49 666 51
rect 660 47 666 49
rect 679 51 685 53
rect 700 55 707 57
rect 700 53 702 55
rect 704 53 707 55
rect 679 49 681 51
rect 683 49 685 51
rect 679 47 685 49
rect 660 43 664 47
rect 651 40 656 43
rect 594 34 599 39
rect 649 38 656 40
rect 649 36 651 38
rect 653 36 656 38
rect 649 34 656 36
rect 658 40 664 43
rect 680 40 685 47
rect 700 47 707 53
rect 784 55 790 57
rect 784 53 786 55
rect 788 53 790 55
rect 784 51 790 53
rect 805 55 812 57
rect 805 53 807 55
rect 809 53 812 55
rect 768 48 773 51
rect 700 45 709 47
rect 658 34 666 40
rect 668 38 676 40
rect 668 36 671 38
rect 673 36 676 38
rect 668 34 676 36
rect 678 34 685 40
rect 689 43 696 45
rect 689 41 691 43
rect 693 41 696 43
rect 689 39 696 41
rect 691 36 696 39
rect 698 36 709 45
rect 711 36 716 47
rect 718 45 725 47
rect 718 43 721 45
rect 723 43 725 45
rect 744 46 753 48
rect 744 44 746 46
rect 748 44 753 46
rect 744 43 753 44
rect 718 41 725 43
rect 718 36 723 41
rect 732 40 737 43
rect 730 38 737 40
rect 730 36 732 38
rect 734 36 737 38
rect 730 34 737 36
rect 739 39 753 43
rect 755 43 763 48
rect 755 41 758 43
rect 760 41 763 43
rect 755 39 763 41
rect 765 45 773 48
rect 765 43 768 45
rect 770 43 773 45
rect 765 39 773 43
rect 775 39 780 51
rect 782 39 790 51
rect 805 47 812 53
rect 889 55 895 57
rect 889 53 891 55
rect 893 53 895 55
rect 889 51 895 53
rect 910 51 916 53
rect 873 48 878 51
rect 805 45 814 47
rect 794 43 801 45
rect 794 41 796 43
rect 798 41 801 43
rect 794 39 801 41
rect 739 34 744 39
rect 796 36 801 39
rect 803 36 814 45
rect 816 36 821 47
rect 823 45 830 47
rect 823 43 826 45
rect 828 43 830 45
rect 849 46 858 48
rect 849 44 851 46
rect 853 44 858 46
rect 849 43 858 44
rect 823 41 830 43
rect 823 36 828 41
rect 837 40 842 43
rect 835 38 842 40
rect 835 36 837 38
rect 839 36 842 38
rect 835 34 842 36
rect 844 39 858 43
rect 860 43 868 48
rect 860 41 863 43
rect 865 41 868 43
rect 860 39 868 41
rect 870 45 878 48
rect 870 43 873 45
rect 875 43 878 45
rect 870 39 878 43
rect 880 39 885 51
rect 887 39 895 51
rect 910 49 912 51
rect 914 49 916 51
rect 910 47 916 49
rect 929 51 935 53
rect 950 55 957 57
rect 950 53 952 55
rect 954 53 957 55
rect 929 49 931 51
rect 933 49 935 51
rect 929 47 935 49
rect 910 43 914 47
rect 901 40 906 43
rect 844 34 849 39
rect 899 38 906 40
rect 899 36 901 38
rect 903 36 906 38
rect 899 34 906 36
rect 908 40 914 43
rect 930 40 935 47
rect 950 47 957 53
rect 1034 55 1040 57
rect 1034 53 1036 55
rect 1038 53 1040 55
rect 1034 51 1040 53
rect 1055 55 1062 57
rect 1055 53 1057 55
rect 1059 53 1062 55
rect 1018 48 1023 51
rect 950 45 959 47
rect 908 34 916 40
rect 918 38 926 40
rect 918 36 921 38
rect 923 36 926 38
rect 918 34 926 36
rect 928 34 935 40
rect 939 43 946 45
rect 939 41 941 43
rect 943 41 946 43
rect 939 39 946 41
rect 941 36 946 39
rect 948 36 959 45
rect 961 36 966 47
rect 968 45 975 47
rect 968 43 971 45
rect 973 43 975 45
rect 994 46 1003 48
rect 994 44 996 46
rect 998 44 1003 46
rect 994 43 1003 44
rect 968 41 975 43
rect 968 36 973 41
rect 982 40 987 43
rect 980 38 987 40
rect 980 36 982 38
rect 984 36 987 38
rect 980 34 987 36
rect 989 39 1003 43
rect 1005 43 1013 48
rect 1005 41 1008 43
rect 1010 41 1013 43
rect 1005 39 1013 41
rect 1015 45 1023 48
rect 1015 43 1018 45
rect 1020 43 1023 45
rect 1015 39 1023 43
rect 1025 39 1030 51
rect 1032 39 1040 51
rect 1055 47 1062 53
rect 1139 55 1145 57
rect 1139 53 1141 55
rect 1143 53 1145 55
rect 1139 51 1145 53
rect 1123 48 1128 51
rect 1055 45 1064 47
rect 1044 43 1051 45
rect 1044 41 1046 43
rect 1048 41 1051 43
rect 1044 39 1051 41
rect 989 34 994 39
rect 1046 36 1051 39
rect 1053 36 1064 45
rect 1066 36 1071 47
rect 1073 45 1080 47
rect 1073 43 1076 45
rect 1078 43 1080 45
rect 1099 46 1108 48
rect 1099 44 1101 46
rect 1103 44 1108 46
rect 1099 43 1108 44
rect 1073 41 1080 43
rect 1073 36 1078 41
rect 1087 40 1092 43
rect 1085 38 1092 40
rect 1085 36 1087 38
rect 1089 36 1092 38
rect 1085 34 1092 36
rect 1094 39 1108 43
rect 1110 43 1118 48
rect 1110 41 1113 43
rect 1115 41 1118 43
rect 1110 39 1118 41
rect 1120 45 1128 48
rect 1120 43 1123 45
rect 1125 43 1128 45
rect 1120 39 1128 43
rect 1130 39 1135 51
rect 1137 39 1145 51
rect 1094 34 1099 39
<< pdif >>
rect 222 302 228 309
rect 201 293 208 302
rect 201 291 203 293
rect 205 291 208 293
rect 201 289 208 291
rect 210 300 218 302
rect 210 298 213 300
rect 215 298 218 300
rect 210 293 218 298
rect 210 291 213 293
rect 215 291 218 293
rect 210 289 218 291
rect 220 295 228 302
rect 220 293 223 295
rect 225 293 228 295
rect 220 291 228 293
rect 230 307 237 309
rect 230 305 233 307
rect 235 305 237 307
rect 230 300 237 305
rect 262 302 268 309
rect 230 298 233 300
rect 235 298 237 300
rect 230 296 237 298
rect 230 291 235 296
rect 241 293 248 302
rect 241 291 243 293
rect 245 291 248 293
rect 220 289 226 291
rect 241 289 248 291
rect 250 300 258 302
rect 250 298 253 300
rect 255 298 258 300
rect 250 293 258 298
rect 250 291 253 293
rect 255 291 258 293
rect 250 289 258 291
rect 260 295 268 302
rect 260 293 263 295
rect 265 293 268 295
rect 260 291 268 293
rect 270 307 277 309
rect 270 305 273 307
rect 275 305 277 307
rect 270 300 277 305
rect 270 298 273 300
rect 275 298 277 300
rect 270 296 277 298
rect 270 291 275 296
rect 290 294 295 309
rect 288 292 295 294
rect 260 289 266 291
rect 288 290 290 292
rect 292 290 295 292
rect 288 288 295 290
rect 290 282 295 288
rect 297 300 305 309
rect 297 298 300 300
rect 302 298 305 300
rect 297 291 305 298
rect 307 307 315 309
rect 307 305 310 307
rect 312 305 315 307
rect 307 300 315 305
rect 307 298 310 300
rect 312 298 315 300
rect 307 291 315 298
rect 317 293 331 309
rect 317 291 326 293
rect 328 291 331 293
rect 297 282 302 291
rect 319 286 331 291
rect 319 284 326 286
rect 328 284 331 286
rect 319 282 331 284
rect 333 307 340 309
rect 333 305 336 307
rect 338 305 340 307
rect 333 303 340 305
rect 333 282 338 303
rect 374 302 380 309
rect 353 293 360 302
rect 353 291 355 293
rect 357 291 360 293
rect 353 289 360 291
rect 362 300 370 302
rect 362 298 365 300
rect 367 298 370 300
rect 362 293 370 298
rect 362 291 365 293
rect 367 291 370 293
rect 362 289 370 291
rect 372 295 380 302
rect 372 293 375 295
rect 377 293 380 295
rect 372 291 380 293
rect 382 307 389 309
rect 382 305 385 307
rect 387 305 389 307
rect 382 300 389 305
rect 438 302 444 309
rect 382 298 385 300
rect 387 298 389 300
rect 382 296 389 298
rect 382 291 387 296
rect 417 293 424 302
rect 417 291 419 293
rect 421 291 424 293
rect 372 289 378 291
rect 417 289 424 291
rect 426 300 434 302
rect 426 298 429 300
rect 431 298 434 300
rect 426 293 434 298
rect 426 291 429 293
rect 431 291 434 293
rect 426 289 434 291
rect 436 295 444 302
rect 436 293 439 295
rect 441 293 444 295
rect 436 291 444 293
rect 446 307 453 309
rect 446 305 449 307
rect 451 305 453 307
rect 446 300 453 305
rect 478 302 484 309
rect 446 298 449 300
rect 451 298 453 300
rect 446 296 453 298
rect 446 291 451 296
rect 457 293 464 302
rect 457 291 459 293
rect 461 291 464 293
rect 436 289 442 291
rect 457 289 464 291
rect 466 300 474 302
rect 466 298 469 300
rect 471 298 474 300
rect 466 293 474 298
rect 466 291 469 293
rect 471 291 474 293
rect 466 289 474 291
rect 476 295 484 302
rect 476 293 479 295
rect 481 293 484 295
rect 476 291 484 293
rect 486 307 493 309
rect 486 305 489 307
rect 491 305 493 307
rect 486 300 493 305
rect 486 298 489 300
rect 491 298 493 300
rect 486 296 493 298
rect 486 291 491 296
rect 506 294 511 309
rect 504 292 511 294
rect 476 289 482 291
rect 504 290 506 292
rect 508 290 511 292
rect 504 288 511 290
rect 506 282 511 288
rect 513 300 521 309
rect 513 298 516 300
rect 518 298 521 300
rect 513 291 521 298
rect 523 307 531 309
rect 523 305 526 307
rect 528 305 531 307
rect 523 300 531 305
rect 523 298 526 300
rect 528 298 531 300
rect 523 291 531 298
rect 533 293 547 309
rect 533 291 542 293
rect 544 291 547 293
rect 513 282 518 291
rect 535 286 547 291
rect 535 284 542 286
rect 544 284 547 286
rect 535 282 547 284
rect 549 307 556 309
rect 549 305 552 307
rect 554 305 556 307
rect 549 303 556 305
rect 549 282 554 303
rect 590 302 596 309
rect 569 293 576 302
rect 569 291 571 293
rect 573 291 576 293
rect 569 289 576 291
rect 578 300 586 302
rect 578 298 581 300
rect 583 298 586 300
rect 578 293 586 298
rect 578 291 581 293
rect 583 291 586 293
rect 578 289 586 291
rect 588 295 596 302
rect 588 293 591 295
rect 593 293 596 295
rect 588 291 596 293
rect 598 307 605 309
rect 598 305 601 307
rect 603 305 605 307
rect 598 300 605 305
rect 643 302 649 309
rect 598 298 601 300
rect 603 298 605 300
rect 598 296 605 298
rect 598 291 603 296
rect 622 293 629 302
rect 622 291 624 293
rect 626 291 629 293
rect 588 289 594 291
rect 622 289 629 291
rect 631 300 639 302
rect 631 298 634 300
rect 636 298 639 300
rect 631 293 639 298
rect 631 291 634 293
rect 636 291 639 293
rect 631 289 639 291
rect 641 295 649 302
rect 641 293 644 295
rect 646 293 649 295
rect 641 291 649 293
rect 651 307 658 309
rect 651 305 654 307
rect 656 305 658 307
rect 651 300 658 305
rect 683 302 689 309
rect 651 298 654 300
rect 656 298 658 300
rect 651 296 658 298
rect 651 291 656 296
rect 662 293 669 302
rect 662 291 664 293
rect 666 291 669 293
rect 641 289 647 291
rect 662 289 669 291
rect 671 300 679 302
rect 671 298 674 300
rect 676 298 679 300
rect 671 293 679 298
rect 671 291 674 293
rect 676 291 679 293
rect 671 289 679 291
rect 681 295 689 302
rect 681 293 684 295
rect 686 293 689 295
rect 681 291 689 293
rect 691 307 698 309
rect 691 305 694 307
rect 696 305 698 307
rect 691 300 698 305
rect 691 298 694 300
rect 696 298 698 300
rect 691 296 698 298
rect 691 291 696 296
rect 711 294 716 309
rect 709 292 716 294
rect 681 289 687 291
rect 709 290 711 292
rect 713 290 716 292
rect 709 288 716 290
rect 711 282 716 288
rect 718 300 726 309
rect 718 298 721 300
rect 723 298 726 300
rect 718 291 726 298
rect 728 307 736 309
rect 728 305 731 307
rect 733 305 736 307
rect 728 300 736 305
rect 728 298 731 300
rect 733 298 736 300
rect 728 291 736 298
rect 738 293 752 309
rect 738 291 747 293
rect 749 291 752 293
rect 718 282 723 291
rect 740 286 752 291
rect 740 284 747 286
rect 749 284 752 286
rect 740 282 752 284
rect 754 307 761 309
rect 754 305 757 307
rect 759 305 761 307
rect 754 303 761 305
rect 754 282 759 303
rect 795 302 801 309
rect 774 293 781 302
rect 774 291 776 293
rect 778 291 781 293
rect 774 289 781 291
rect 783 300 791 302
rect 783 298 786 300
rect 788 298 791 300
rect 783 293 791 298
rect 783 291 786 293
rect 788 291 791 293
rect 783 289 791 291
rect 793 295 801 302
rect 793 293 796 295
rect 798 293 801 295
rect 793 291 801 293
rect 803 307 810 309
rect 803 305 806 307
rect 808 305 810 307
rect 803 300 810 305
rect 862 302 868 309
rect 803 298 806 300
rect 808 298 810 300
rect 803 296 810 298
rect 803 291 808 296
rect 841 293 848 302
rect 841 291 843 293
rect 845 291 848 293
rect 793 289 799 291
rect 841 289 848 291
rect 850 300 858 302
rect 850 298 853 300
rect 855 298 858 300
rect 850 293 858 298
rect 850 291 853 293
rect 855 291 858 293
rect 850 289 858 291
rect 860 295 868 302
rect 860 293 863 295
rect 865 293 868 295
rect 860 291 868 293
rect 870 307 877 309
rect 870 305 873 307
rect 875 305 877 307
rect 870 300 877 305
rect 902 302 908 309
rect 870 298 873 300
rect 875 298 877 300
rect 870 296 877 298
rect 870 291 875 296
rect 881 293 888 302
rect 881 291 883 293
rect 885 291 888 293
rect 860 289 866 291
rect 881 289 888 291
rect 890 300 898 302
rect 890 298 893 300
rect 895 298 898 300
rect 890 293 898 298
rect 890 291 893 293
rect 895 291 898 293
rect 890 289 898 291
rect 900 295 908 302
rect 900 293 903 295
rect 905 293 908 295
rect 900 291 908 293
rect 910 307 917 309
rect 910 305 913 307
rect 915 305 917 307
rect 910 300 917 305
rect 910 298 913 300
rect 915 298 917 300
rect 910 296 917 298
rect 910 291 915 296
rect 930 294 935 309
rect 928 292 935 294
rect 900 289 906 291
rect 928 290 930 292
rect 932 290 935 292
rect 928 288 935 290
rect 930 282 935 288
rect 937 300 945 309
rect 937 298 940 300
rect 942 298 945 300
rect 937 291 945 298
rect 947 307 955 309
rect 947 305 950 307
rect 952 305 955 307
rect 947 300 955 305
rect 947 298 950 300
rect 952 298 955 300
rect 947 291 955 298
rect 957 293 971 309
rect 957 291 966 293
rect 968 291 971 293
rect 937 282 942 291
rect 959 286 971 291
rect 959 284 966 286
rect 968 284 971 286
rect 959 282 971 284
rect 973 307 980 309
rect 973 305 976 307
rect 978 305 980 307
rect 973 303 980 305
rect 973 282 978 303
rect 1014 302 1020 309
rect 993 293 1000 302
rect 993 291 995 293
rect 997 291 1000 293
rect 993 289 1000 291
rect 1002 300 1010 302
rect 1002 298 1005 300
rect 1007 298 1010 300
rect 1002 293 1010 298
rect 1002 291 1005 293
rect 1007 291 1010 293
rect 1002 289 1010 291
rect 1012 295 1020 302
rect 1012 293 1015 295
rect 1017 293 1020 295
rect 1012 291 1020 293
rect 1022 307 1029 309
rect 1022 305 1025 307
rect 1027 305 1029 307
rect 1022 300 1029 305
rect 1022 298 1025 300
rect 1027 298 1029 300
rect 1022 296 1029 298
rect 1022 291 1027 296
rect 1012 289 1018 291
rect 212 261 218 263
rect 203 256 208 261
rect 201 254 208 256
rect 201 252 203 254
rect 205 252 208 254
rect 201 247 208 252
rect 201 245 203 247
rect 205 245 208 247
rect 201 243 208 245
rect 210 259 218 261
rect 210 257 213 259
rect 215 257 218 259
rect 210 250 218 257
rect 220 261 228 263
rect 220 259 223 261
rect 225 259 228 261
rect 220 254 228 259
rect 220 252 223 254
rect 225 252 228 254
rect 220 250 228 252
rect 230 261 237 263
rect 230 259 233 261
rect 235 259 237 261
rect 230 250 237 259
rect 241 261 248 263
rect 241 259 243 261
rect 245 259 248 261
rect 241 250 248 259
rect 250 261 258 263
rect 250 259 253 261
rect 255 259 258 261
rect 250 254 258 259
rect 250 252 253 254
rect 255 252 258 254
rect 250 250 258 252
rect 260 261 266 263
rect 292 261 298 263
rect 260 259 268 261
rect 260 257 263 259
rect 265 257 268 259
rect 260 250 268 257
rect 210 243 216 250
rect 262 243 268 250
rect 270 256 275 261
rect 283 256 288 261
rect 270 254 277 256
rect 270 252 273 254
rect 275 252 277 254
rect 270 247 277 252
rect 270 245 273 247
rect 275 245 277 247
rect 270 243 277 245
rect 281 254 288 256
rect 281 252 283 254
rect 285 252 288 254
rect 281 247 288 252
rect 281 245 283 247
rect 285 245 288 247
rect 281 243 288 245
rect 290 259 298 261
rect 290 257 293 259
rect 295 257 298 259
rect 290 250 298 257
rect 300 261 308 263
rect 300 259 303 261
rect 305 259 308 261
rect 300 254 308 259
rect 300 252 303 254
rect 305 252 308 254
rect 300 250 308 252
rect 310 261 317 263
rect 310 259 313 261
rect 315 259 317 261
rect 310 250 317 259
rect 290 243 296 250
rect 332 249 337 270
rect 330 247 337 249
rect 330 245 332 247
rect 334 245 337 247
rect 330 243 337 245
rect 339 268 351 270
rect 339 266 342 268
rect 344 266 351 268
rect 339 261 351 266
rect 368 261 373 270
rect 339 259 342 261
rect 344 259 353 261
rect 339 243 353 259
rect 355 254 363 261
rect 355 252 358 254
rect 360 252 363 254
rect 355 247 363 252
rect 355 245 358 247
rect 360 245 363 247
rect 355 243 363 245
rect 365 254 373 261
rect 365 252 368 254
rect 370 252 373 254
rect 365 243 373 252
rect 375 264 380 270
rect 375 262 382 264
rect 375 260 378 262
rect 380 260 382 262
rect 428 261 434 263
rect 375 258 382 260
rect 375 243 380 258
rect 419 256 424 261
rect 417 254 424 256
rect 417 252 419 254
rect 421 252 424 254
rect 417 247 424 252
rect 417 245 419 247
rect 421 245 424 247
rect 417 243 424 245
rect 426 259 434 261
rect 426 257 429 259
rect 431 257 434 259
rect 426 250 434 257
rect 436 261 444 263
rect 436 259 439 261
rect 441 259 444 261
rect 436 254 444 259
rect 436 252 439 254
rect 441 252 444 254
rect 436 250 444 252
rect 446 261 453 263
rect 446 259 449 261
rect 451 259 453 261
rect 446 250 453 259
rect 457 261 464 263
rect 457 259 459 261
rect 461 259 464 261
rect 457 250 464 259
rect 466 261 474 263
rect 466 259 469 261
rect 471 259 474 261
rect 466 254 474 259
rect 466 252 469 254
rect 471 252 474 254
rect 466 250 474 252
rect 476 261 482 263
rect 508 261 514 263
rect 476 259 484 261
rect 476 257 479 259
rect 481 257 484 259
rect 476 250 484 257
rect 426 243 432 250
rect 478 243 484 250
rect 486 256 491 261
rect 499 256 504 261
rect 486 254 493 256
rect 486 252 489 254
rect 491 252 493 254
rect 486 247 493 252
rect 486 245 489 247
rect 491 245 493 247
rect 486 243 493 245
rect 497 254 504 256
rect 497 252 499 254
rect 501 252 504 254
rect 497 247 504 252
rect 497 245 499 247
rect 501 245 504 247
rect 497 243 504 245
rect 506 259 514 261
rect 506 257 509 259
rect 511 257 514 259
rect 506 250 514 257
rect 516 261 524 263
rect 516 259 519 261
rect 521 259 524 261
rect 516 254 524 259
rect 516 252 519 254
rect 521 252 524 254
rect 516 250 524 252
rect 526 261 533 263
rect 526 259 529 261
rect 531 259 533 261
rect 526 250 533 259
rect 506 243 512 250
rect 548 249 553 270
rect 546 247 553 249
rect 546 245 548 247
rect 550 245 553 247
rect 546 243 553 245
rect 555 268 567 270
rect 555 266 558 268
rect 560 266 567 268
rect 555 261 567 266
rect 584 261 589 270
rect 555 259 558 261
rect 560 259 569 261
rect 555 243 569 259
rect 571 254 579 261
rect 571 252 574 254
rect 576 252 579 254
rect 571 247 579 252
rect 571 245 574 247
rect 576 245 579 247
rect 571 243 579 245
rect 581 254 589 261
rect 581 252 584 254
rect 586 252 589 254
rect 581 243 589 252
rect 591 264 596 270
rect 591 262 598 264
rect 591 260 594 262
rect 596 260 598 262
rect 633 261 639 263
rect 591 258 598 260
rect 591 243 596 258
rect 624 256 629 261
rect 622 254 629 256
rect 622 252 624 254
rect 626 252 629 254
rect 622 247 629 252
rect 622 245 624 247
rect 626 245 629 247
rect 622 243 629 245
rect 631 259 639 261
rect 631 257 634 259
rect 636 257 639 259
rect 631 250 639 257
rect 641 261 649 263
rect 641 259 644 261
rect 646 259 649 261
rect 641 254 649 259
rect 641 252 644 254
rect 646 252 649 254
rect 641 250 649 252
rect 651 261 658 263
rect 651 259 654 261
rect 656 259 658 261
rect 651 250 658 259
rect 662 261 669 263
rect 662 259 664 261
rect 666 259 669 261
rect 662 250 669 259
rect 671 261 679 263
rect 671 259 674 261
rect 676 259 679 261
rect 671 254 679 259
rect 671 252 674 254
rect 676 252 679 254
rect 671 250 679 252
rect 681 261 687 263
rect 713 261 719 263
rect 681 259 689 261
rect 681 257 684 259
rect 686 257 689 259
rect 681 250 689 257
rect 631 243 637 250
rect 683 243 689 250
rect 691 256 696 261
rect 704 256 709 261
rect 691 254 698 256
rect 691 252 694 254
rect 696 252 698 254
rect 691 247 698 252
rect 691 245 694 247
rect 696 245 698 247
rect 691 243 698 245
rect 702 254 709 256
rect 702 252 704 254
rect 706 252 709 254
rect 702 247 709 252
rect 702 245 704 247
rect 706 245 709 247
rect 702 243 709 245
rect 711 259 719 261
rect 711 257 714 259
rect 716 257 719 259
rect 711 250 719 257
rect 721 261 729 263
rect 721 259 724 261
rect 726 259 729 261
rect 721 254 729 259
rect 721 252 724 254
rect 726 252 729 254
rect 721 250 729 252
rect 731 261 738 263
rect 731 259 734 261
rect 736 259 738 261
rect 731 250 738 259
rect 711 243 717 250
rect 753 249 758 270
rect 751 247 758 249
rect 751 245 753 247
rect 755 245 758 247
rect 751 243 758 245
rect 760 268 772 270
rect 760 266 763 268
rect 765 266 772 268
rect 760 261 772 266
rect 789 261 794 270
rect 760 259 763 261
rect 765 259 774 261
rect 760 243 774 259
rect 776 254 784 261
rect 776 252 779 254
rect 781 252 784 254
rect 776 247 784 252
rect 776 245 779 247
rect 781 245 784 247
rect 776 243 784 245
rect 786 254 794 261
rect 786 252 789 254
rect 791 252 794 254
rect 786 243 794 252
rect 796 264 801 270
rect 796 262 803 264
rect 796 260 799 262
rect 801 260 803 262
rect 852 261 858 263
rect 796 258 803 260
rect 796 243 801 258
rect 843 256 848 261
rect 841 254 848 256
rect 841 252 843 254
rect 845 252 848 254
rect 841 247 848 252
rect 841 245 843 247
rect 845 245 848 247
rect 841 243 848 245
rect 850 259 858 261
rect 850 257 853 259
rect 855 257 858 259
rect 850 250 858 257
rect 860 261 868 263
rect 860 259 863 261
rect 865 259 868 261
rect 860 254 868 259
rect 860 252 863 254
rect 865 252 868 254
rect 860 250 868 252
rect 870 261 877 263
rect 870 259 873 261
rect 875 259 877 261
rect 870 250 877 259
rect 881 261 888 263
rect 881 259 883 261
rect 885 259 888 261
rect 881 250 888 259
rect 890 261 898 263
rect 890 259 893 261
rect 895 259 898 261
rect 890 254 898 259
rect 890 252 893 254
rect 895 252 898 254
rect 890 250 898 252
rect 900 261 906 263
rect 932 261 938 263
rect 900 259 908 261
rect 900 257 903 259
rect 905 257 908 259
rect 900 250 908 257
rect 850 243 856 250
rect 902 243 908 250
rect 910 256 915 261
rect 923 256 928 261
rect 910 254 917 256
rect 910 252 913 254
rect 915 252 917 254
rect 910 247 917 252
rect 910 245 913 247
rect 915 245 917 247
rect 910 243 917 245
rect 921 254 928 256
rect 921 252 923 254
rect 925 252 928 254
rect 921 247 928 252
rect 921 245 923 247
rect 925 245 928 247
rect 921 243 928 245
rect 930 259 938 261
rect 930 257 933 259
rect 935 257 938 259
rect 930 250 938 257
rect 940 261 948 263
rect 940 259 943 261
rect 945 259 948 261
rect 940 254 948 259
rect 940 252 943 254
rect 945 252 948 254
rect 940 250 948 252
rect 950 261 957 263
rect 950 259 953 261
rect 955 259 957 261
rect 950 250 957 259
rect 930 243 936 250
rect 972 249 977 270
rect 970 247 977 249
rect 970 245 972 247
rect 974 245 977 247
rect 970 243 977 245
rect 979 268 991 270
rect 979 266 982 268
rect 984 266 991 268
rect 979 261 991 266
rect 1008 261 1013 270
rect 979 259 982 261
rect 984 259 993 261
rect 979 243 993 259
rect 995 254 1003 261
rect 995 252 998 254
rect 1000 252 1003 254
rect 995 247 1003 252
rect 995 245 998 247
rect 1000 245 1003 247
rect 995 243 1003 245
rect 1005 254 1013 261
rect 1005 252 1008 254
rect 1010 252 1013 254
rect 1005 243 1013 252
rect 1015 264 1020 270
rect 1015 262 1022 264
rect 1015 260 1018 262
rect 1020 260 1022 262
rect 1056 261 1062 263
rect 1015 258 1022 260
rect 1015 243 1020 258
rect 1047 256 1052 261
rect 1045 254 1052 256
rect 1045 252 1047 254
rect 1049 252 1052 254
rect 1045 247 1052 252
rect 1045 245 1047 247
rect 1049 245 1052 247
rect 1045 243 1052 245
rect 1054 259 1062 261
rect 1054 257 1057 259
rect 1059 257 1062 259
rect 1054 250 1062 257
rect 1064 261 1072 263
rect 1064 259 1067 261
rect 1069 259 1072 261
rect 1064 254 1072 259
rect 1064 252 1067 254
rect 1069 252 1072 254
rect 1064 250 1072 252
rect 1074 261 1081 263
rect 1074 259 1077 261
rect 1079 259 1081 261
rect 1074 250 1081 259
rect 1054 243 1060 250
rect 1096 249 1101 270
rect 1094 247 1101 249
rect 1094 245 1096 247
rect 1098 245 1101 247
rect 1094 243 1101 245
rect 1103 268 1115 270
rect 1103 266 1106 268
rect 1108 266 1115 268
rect 1103 261 1115 266
rect 1132 261 1137 270
rect 1103 259 1106 261
rect 1108 259 1117 261
rect 1103 243 1117 259
rect 1119 254 1127 261
rect 1119 252 1122 254
rect 1124 252 1127 254
rect 1119 247 1127 252
rect 1119 245 1122 247
rect 1124 245 1127 247
rect 1119 243 1127 245
rect 1129 254 1137 261
rect 1129 252 1132 254
rect 1134 252 1137 254
rect 1129 243 1137 252
rect 1139 264 1144 270
rect 1139 262 1146 264
rect 1139 260 1142 262
rect 1144 260 1146 262
rect 1139 258 1146 260
rect 1139 243 1144 258
rect 153 161 158 166
rect 151 159 158 161
rect 151 157 153 159
rect 155 157 158 159
rect 151 152 158 157
rect 151 150 153 152
rect 155 150 158 152
rect 151 148 158 150
rect 160 159 168 166
rect 191 163 198 165
rect 191 161 193 163
rect 195 161 198 163
rect 160 148 171 159
rect 162 142 171 148
rect 162 140 164 142
rect 166 140 171 142
rect 162 138 171 140
rect 173 138 178 159
rect 180 151 185 159
rect 191 156 198 161
rect 191 154 193 156
rect 195 154 198 156
rect 191 152 198 154
rect 180 149 187 151
rect 180 147 183 149
rect 185 147 187 149
rect 193 147 198 152
rect 200 158 206 165
rect 240 163 247 165
rect 240 161 242 163
rect 244 161 247 163
rect 240 159 247 161
rect 200 151 208 158
rect 200 149 203 151
rect 205 149 208 151
rect 200 147 208 149
rect 180 145 187 147
rect 180 138 185 145
rect 202 145 208 147
rect 210 156 218 158
rect 210 154 213 156
rect 215 154 218 156
rect 210 149 218 154
rect 210 147 213 149
rect 215 147 218 149
rect 210 145 218 147
rect 220 149 227 158
rect 220 147 223 149
rect 225 147 227 149
rect 220 145 227 147
rect 242 138 247 159
rect 249 149 263 165
rect 249 147 252 149
rect 254 147 263 149
rect 265 163 273 165
rect 265 161 268 163
rect 270 161 273 163
rect 265 156 273 161
rect 265 154 268 156
rect 270 154 273 156
rect 265 147 273 154
rect 275 156 283 165
rect 275 154 278 156
rect 280 154 283 156
rect 275 147 283 154
rect 249 142 261 147
rect 249 140 252 142
rect 254 140 261 142
rect 249 138 261 140
rect 278 138 283 147
rect 285 150 290 165
rect 296 163 303 165
rect 296 161 298 163
rect 300 161 303 163
rect 296 156 303 161
rect 296 154 298 156
rect 300 154 303 156
rect 296 152 303 154
rect 285 148 292 150
rect 285 146 288 148
rect 290 146 292 148
rect 298 147 303 152
rect 305 158 311 165
rect 345 163 352 165
rect 345 161 347 163
rect 349 161 352 163
rect 345 159 352 161
rect 305 151 313 158
rect 305 149 308 151
rect 310 149 313 151
rect 305 147 313 149
rect 285 144 292 146
rect 285 138 290 144
rect 307 145 313 147
rect 315 156 323 158
rect 315 154 318 156
rect 320 154 323 156
rect 315 149 323 154
rect 315 147 318 149
rect 320 147 323 149
rect 315 145 323 147
rect 325 149 332 158
rect 325 147 328 149
rect 330 147 332 149
rect 325 145 332 147
rect 347 138 352 159
rect 354 149 368 165
rect 354 147 357 149
rect 359 147 368 149
rect 370 163 378 165
rect 370 161 373 163
rect 375 161 378 163
rect 370 156 378 161
rect 370 154 373 156
rect 375 154 378 156
rect 370 147 378 154
rect 380 156 388 165
rect 380 154 383 156
rect 385 154 388 156
rect 380 147 388 154
rect 354 142 366 147
rect 354 140 357 142
rect 359 140 366 142
rect 354 138 366 140
rect 383 138 388 147
rect 390 150 395 165
rect 403 161 408 166
rect 401 159 408 161
rect 401 157 403 159
rect 405 157 408 159
rect 401 152 408 157
rect 401 150 403 152
rect 405 150 408 152
rect 390 148 397 150
rect 401 148 408 150
rect 410 159 418 166
rect 441 163 448 165
rect 441 161 443 163
rect 445 161 448 163
rect 410 148 421 159
rect 390 146 393 148
rect 395 146 397 148
rect 390 144 397 146
rect 390 138 395 144
rect 412 142 421 148
rect 412 140 414 142
rect 416 140 421 142
rect 412 138 421 140
rect 423 138 428 159
rect 430 151 435 159
rect 441 156 448 161
rect 441 154 443 156
rect 445 154 448 156
rect 441 152 448 154
rect 430 149 437 151
rect 430 147 433 149
rect 435 147 437 149
rect 443 147 448 152
rect 450 158 456 165
rect 490 163 497 165
rect 490 161 492 163
rect 494 161 497 163
rect 490 159 497 161
rect 450 151 458 158
rect 450 149 453 151
rect 455 149 458 151
rect 450 147 458 149
rect 430 145 437 147
rect 430 138 435 145
rect 452 145 458 147
rect 460 156 468 158
rect 460 154 463 156
rect 465 154 468 156
rect 460 149 468 154
rect 460 147 463 149
rect 465 147 468 149
rect 460 145 468 147
rect 470 149 477 158
rect 470 147 473 149
rect 475 147 477 149
rect 470 145 477 147
rect 492 138 497 159
rect 499 149 513 165
rect 499 147 502 149
rect 504 147 513 149
rect 515 163 523 165
rect 515 161 518 163
rect 520 161 523 163
rect 515 156 523 161
rect 515 154 518 156
rect 520 154 523 156
rect 515 147 523 154
rect 525 156 533 165
rect 525 154 528 156
rect 530 154 533 156
rect 525 147 533 154
rect 499 142 511 147
rect 499 140 502 142
rect 504 140 511 142
rect 499 138 511 140
rect 528 138 533 147
rect 535 150 540 165
rect 546 163 553 165
rect 546 161 548 163
rect 550 161 553 163
rect 546 156 553 161
rect 546 154 548 156
rect 550 154 553 156
rect 546 152 553 154
rect 535 148 542 150
rect 535 146 538 148
rect 540 146 542 148
rect 548 147 553 152
rect 555 158 561 165
rect 595 163 602 165
rect 595 161 597 163
rect 599 161 602 163
rect 595 159 602 161
rect 555 151 563 158
rect 555 149 558 151
rect 560 149 563 151
rect 555 147 563 149
rect 535 144 542 146
rect 535 138 540 144
rect 557 145 563 147
rect 565 156 573 158
rect 565 154 568 156
rect 570 154 573 156
rect 565 149 573 154
rect 565 147 568 149
rect 570 147 573 149
rect 565 145 573 147
rect 575 149 582 158
rect 575 147 578 149
rect 580 147 582 149
rect 575 145 582 147
rect 597 138 602 159
rect 604 149 618 165
rect 604 147 607 149
rect 609 147 618 149
rect 620 163 628 165
rect 620 161 623 163
rect 625 161 628 163
rect 620 156 628 161
rect 620 154 623 156
rect 625 154 628 156
rect 620 147 628 154
rect 630 156 638 165
rect 630 154 633 156
rect 635 154 638 156
rect 630 147 638 154
rect 604 142 616 147
rect 604 140 607 142
rect 609 140 616 142
rect 604 138 616 140
rect 633 138 638 147
rect 640 150 645 165
rect 653 161 658 166
rect 651 159 658 161
rect 651 157 653 159
rect 655 157 658 159
rect 651 152 658 157
rect 651 150 653 152
rect 655 150 658 152
rect 640 148 647 150
rect 651 148 658 150
rect 660 159 668 166
rect 691 163 698 165
rect 691 161 693 163
rect 695 161 698 163
rect 660 148 671 159
rect 640 146 643 148
rect 645 146 647 148
rect 640 144 647 146
rect 640 138 645 144
rect 662 142 671 148
rect 662 140 664 142
rect 666 140 671 142
rect 662 138 671 140
rect 673 138 678 159
rect 680 151 685 159
rect 691 156 698 161
rect 691 154 693 156
rect 695 154 698 156
rect 691 152 698 154
rect 680 149 687 151
rect 680 147 683 149
rect 685 147 687 149
rect 693 147 698 152
rect 700 158 706 165
rect 740 163 747 165
rect 740 161 742 163
rect 744 161 747 163
rect 740 159 747 161
rect 700 151 708 158
rect 700 149 703 151
rect 705 149 708 151
rect 700 147 708 149
rect 680 145 687 147
rect 680 138 685 145
rect 702 145 708 147
rect 710 156 718 158
rect 710 154 713 156
rect 715 154 718 156
rect 710 149 718 154
rect 710 147 713 149
rect 715 147 718 149
rect 710 145 718 147
rect 720 149 727 158
rect 720 147 723 149
rect 725 147 727 149
rect 720 145 727 147
rect 742 138 747 159
rect 749 149 763 165
rect 749 147 752 149
rect 754 147 763 149
rect 765 163 773 165
rect 765 161 768 163
rect 770 161 773 163
rect 765 156 773 161
rect 765 154 768 156
rect 770 154 773 156
rect 765 147 773 154
rect 775 156 783 165
rect 775 154 778 156
rect 780 154 783 156
rect 775 147 783 154
rect 749 142 761 147
rect 749 140 752 142
rect 754 140 761 142
rect 749 138 761 140
rect 778 138 783 147
rect 785 150 790 165
rect 796 163 803 165
rect 796 161 798 163
rect 800 161 803 163
rect 796 156 803 161
rect 796 154 798 156
rect 800 154 803 156
rect 796 152 803 154
rect 785 148 792 150
rect 785 146 788 148
rect 790 146 792 148
rect 798 147 803 152
rect 805 158 811 165
rect 845 163 852 165
rect 845 161 847 163
rect 849 161 852 163
rect 845 159 852 161
rect 805 151 813 158
rect 805 149 808 151
rect 810 149 813 151
rect 805 147 813 149
rect 785 144 792 146
rect 785 138 790 144
rect 807 145 813 147
rect 815 156 823 158
rect 815 154 818 156
rect 820 154 823 156
rect 815 149 823 154
rect 815 147 818 149
rect 820 147 823 149
rect 815 145 823 147
rect 825 149 832 158
rect 825 147 828 149
rect 830 147 832 149
rect 825 145 832 147
rect 847 138 852 159
rect 854 149 868 165
rect 854 147 857 149
rect 859 147 868 149
rect 870 163 878 165
rect 870 161 873 163
rect 875 161 878 163
rect 870 156 878 161
rect 870 154 873 156
rect 875 154 878 156
rect 870 147 878 154
rect 880 156 888 165
rect 880 154 883 156
rect 885 154 888 156
rect 880 147 888 154
rect 854 142 866 147
rect 854 140 857 142
rect 859 140 866 142
rect 854 138 866 140
rect 883 138 888 147
rect 890 150 895 165
rect 903 161 908 166
rect 901 159 908 161
rect 901 157 903 159
rect 905 157 908 159
rect 901 152 908 157
rect 901 150 903 152
rect 905 150 908 152
rect 890 148 897 150
rect 901 148 908 150
rect 910 159 918 166
rect 941 163 948 165
rect 941 161 943 163
rect 945 161 948 163
rect 910 148 921 159
rect 890 146 893 148
rect 895 146 897 148
rect 890 144 897 146
rect 890 138 895 144
rect 912 142 921 148
rect 912 140 914 142
rect 916 140 921 142
rect 912 138 921 140
rect 923 138 928 159
rect 930 151 935 159
rect 941 156 948 161
rect 941 154 943 156
rect 945 154 948 156
rect 941 152 948 154
rect 930 149 937 151
rect 930 147 933 149
rect 935 147 937 149
rect 943 147 948 152
rect 950 158 956 165
rect 990 163 997 165
rect 990 161 992 163
rect 994 161 997 163
rect 990 159 997 161
rect 950 151 958 158
rect 950 149 953 151
rect 955 149 958 151
rect 950 147 958 149
rect 930 145 937 147
rect 930 138 935 145
rect 952 145 958 147
rect 960 156 968 158
rect 960 154 963 156
rect 965 154 968 156
rect 960 149 968 154
rect 960 147 963 149
rect 965 147 968 149
rect 960 145 968 147
rect 970 149 977 158
rect 970 147 973 149
rect 975 147 977 149
rect 970 145 977 147
rect 992 138 997 159
rect 999 149 1013 165
rect 999 147 1002 149
rect 1004 147 1013 149
rect 1015 163 1023 165
rect 1015 161 1018 163
rect 1020 161 1023 163
rect 1015 156 1023 161
rect 1015 154 1018 156
rect 1020 154 1023 156
rect 1015 147 1023 154
rect 1025 156 1033 165
rect 1025 154 1028 156
rect 1030 154 1033 156
rect 1025 147 1033 154
rect 999 142 1011 147
rect 999 140 1002 142
rect 1004 140 1011 142
rect 999 138 1011 140
rect 1028 138 1033 147
rect 1035 150 1040 165
rect 1046 163 1053 165
rect 1046 161 1048 163
rect 1050 161 1053 163
rect 1046 156 1053 161
rect 1046 154 1048 156
rect 1050 154 1053 156
rect 1046 152 1053 154
rect 1035 148 1042 150
rect 1035 146 1038 148
rect 1040 146 1042 148
rect 1048 147 1053 152
rect 1055 158 1061 165
rect 1095 163 1102 165
rect 1095 161 1097 163
rect 1099 161 1102 163
rect 1095 159 1102 161
rect 1055 151 1063 158
rect 1055 149 1058 151
rect 1060 149 1063 151
rect 1055 147 1063 149
rect 1035 144 1042 146
rect 1035 138 1040 144
rect 1057 145 1063 147
rect 1065 156 1073 158
rect 1065 154 1068 156
rect 1070 154 1073 156
rect 1065 149 1073 154
rect 1065 147 1068 149
rect 1070 147 1073 149
rect 1065 145 1073 147
rect 1075 149 1082 158
rect 1075 147 1078 149
rect 1080 147 1082 149
rect 1075 145 1082 147
rect 1097 138 1102 159
rect 1104 149 1118 165
rect 1104 147 1107 149
rect 1109 147 1118 149
rect 1120 163 1128 165
rect 1120 161 1123 163
rect 1125 161 1128 163
rect 1120 156 1128 161
rect 1120 154 1123 156
rect 1125 154 1128 156
rect 1120 147 1128 154
rect 1130 156 1138 165
rect 1130 154 1133 156
rect 1135 154 1138 156
rect 1130 147 1138 154
rect 1104 142 1116 147
rect 1104 140 1107 142
rect 1109 140 1116 142
rect 1104 138 1116 140
rect 1133 138 1138 147
rect 1140 150 1145 165
rect 1140 148 1147 150
rect 1140 146 1143 148
rect 1145 146 1147 148
rect 1140 144 1147 146
rect 1140 138 1145 144
rect 161 124 170 126
rect 161 122 163 124
rect 165 122 170 124
rect 161 116 170 122
rect 150 114 157 116
rect 150 112 152 114
rect 154 112 157 114
rect 150 107 157 112
rect 150 105 152 107
rect 154 105 157 107
rect 150 103 157 105
rect 152 98 157 103
rect 159 105 170 116
rect 172 105 177 126
rect 179 119 184 126
rect 179 117 186 119
rect 201 117 207 119
rect 179 115 182 117
rect 184 115 186 117
rect 179 113 186 115
rect 179 105 184 113
rect 192 112 197 117
rect 190 110 197 112
rect 190 108 192 110
rect 194 108 197 110
rect 159 98 167 105
rect 190 103 197 108
rect 190 101 192 103
rect 194 101 197 103
rect 190 99 197 101
rect 199 115 207 117
rect 199 113 202 115
rect 204 113 207 115
rect 199 106 207 113
rect 209 117 217 119
rect 209 115 212 117
rect 214 115 217 117
rect 209 110 217 115
rect 209 108 212 110
rect 214 108 217 110
rect 209 106 217 108
rect 219 117 226 119
rect 219 115 222 117
rect 224 115 226 117
rect 219 106 226 115
rect 199 99 205 106
rect 241 105 246 126
rect 239 103 246 105
rect 239 101 241 103
rect 243 101 246 103
rect 239 99 246 101
rect 248 124 260 126
rect 248 122 251 124
rect 253 122 260 124
rect 248 117 260 122
rect 277 117 282 126
rect 248 115 251 117
rect 253 115 262 117
rect 248 99 262 115
rect 264 110 272 117
rect 264 108 267 110
rect 269 108 272 110
rect 264 103 272 108
rect 264 101 267 103
rect 269 101 272 103
rect 264 99 272 101
rect 274 110 282 117
rect 274 108 277 110
rect 279 108 282 110
rect 274 99 282 108
rect 284 120 289 126
rect 284 118 291 120
rect 284 116 287 118
rect 289 116 291 118
rect 306 117 312 119
rect 284 114 291 116
rect 284 99 289 114
rect 297 112 302 117
rect 295 110 302 112
rect 295 108 297 110
rect 299 108 302 110
rect 295 103 302 108
rect 295 101 297 103
rect 299 101 302 103
rect 295 99 302 101
rect 304 115 312 117
rect 304 113 307 115
rect 309 113 312 115
rect 304 106 312 113
rect 314 117 322 119
rect 314 115 317 117
rect 319 115 322 117
rect 314 110 322 115
rect 314 108 317 110
rect 319 108 322 110
rect 314 106 322 108
rect 324 117 331 119
rect 324 115 327 117
rect 329 115 331 117
rect 324 106 331 115
rect 304 99 310 106
rect 346 105 351 126
rect 344 103 351 105
rect 344 101 346 103
rect 348 101 351 103
rect 344 99 351 101
rect 353 124 365 126
rect 353 122 356 124
rect 358 122 365 124
rect 353 117 365 122
rect 382 117 387 126
rect 353 115 356 117
rect 358 115 367 117
rect 353 99 367 115
rect 369 110 377 117
rect 369 108 372 110
rect 374 108 377 110
rect 369 103 377 108
rect 369 101 372 103
rect 374 101 377 103
rect 369 99 377 101
rect 379 110 387 117
rect 379 108 382 110
rect 384 108 387 110
rect 379 99 387 108
rect 389 120 394 126
rect 411 124 420 126
rect 411 122 413 124
rect 415 122 420 124
rect 389 118 396 120
rect 389 116 392 118
rect 394 116 396 118
rect 411 116 420 122
rect 389 114 396 116
rect 400 114 407 116
rect 389 99 394 114
rect 400 112 402 114
rect 404 112 407 114
rect 400 107 407 112
rect 400 105 402 107
rect 404 105 407 107
rect 400 103 407 105
rect 402 98 407 103
rect 409 105 420 116
rect 422 105 427 126
rect 429 119 434 126
rect 429 117 436 119
rect 451 117 457 119
rect 429 115 432 117
rect 434 115 436 117
rect 429 113 436 115
rect 429 105 434 113
rect 442 112 447 117
rect 440 110 447 112
rect 440 108 442 110
rect 444 108 447 110
rect 409 98 417 105
rect 440 103 447 108
rect 440 101 442 103
rect 444 101 447 103
rect 440 99 447 101
rect 449 115 457 117
rect 449 113 452 115
rect 454 113 457 115
rect 449 106 457 113
rect 459 117 467 119
rect 459 115 462 117
rect 464 115 467 117
rect 459 110 467 115
rect 459 108 462 110
rect 464 108 467 110
rect 459 106 467 108
rect 469 117 476 119
rect 469 115 472 117
rect 474 115 476 117
rect 469 106 476 115
rect 449 99 455 106
rect 491 105 496 126
rect 489 103 496 105
rect 489 101 491 103
rect 493 101 496 103
rect 489 99 496 101
rect 498 124 510 126
rect 498 122 501 124
rect 503 122 510 124
rect 498 117 510 122
rect 527 117 532 126
rect 498 115 501 117
rect 503 115 512 117
rect 498 99 512 115
rect 514 110 522 117
rect 514 108 517 110
rect 519 108 522 110
rect 514 103 522 108
rect 514 101 517 103
rect 519 101 522 103
rect 514 99 522 101
rect 524 110 532 117
rect 524 108 527 110
rect 529 108 532 110
rect 524 99 532 108
rect 534 120 539 126
rect 534 118 541 120
rect 534 116 537 118
rect 539 116 541 118
rect 556 117 562 119
rect 534 114 541 116
rect 534 99 539 114
rect 547 112 552 117
rect 545 110 552 112
rect 545 108 547 110
rect 549 108 552 110
rect 545 103 552 108
rect 545 101 547 103
rect 549 101 552 103
rect 545 99 552 101
rect 554 115 562 117
rect 554 113 557 115
rect 559 113 562 115
rect 554 106 562 113
rect 564 117 572 119
rect 564 115 567 117
rect 569 115 572 117
rect 564 110 572 115
rect 564 108 567 110
rect 569 108 572 110
rect 564 106 572 108
rect 574 117 581 119
rect 574 115 577 117
rect 579 115 581 117
rect 574 106 581 115
rect 554 99 560 106
rect 596 105 601 126
rect 594 103 601 105
rect 594 101 596 103
rect 598 101 601 103
rect 594 99 601 101
rect 603 124 615 126
rect 603 122 606 124
rect 608 122 615 124
rect 603 117 615 122
rect 632 117 637 126
rect 603 115 606 117
rect 608 115 617 117
rect 603 99 617 115
rect 619 110 627 117
rect 619 108 622 110
rect 624 108 627 110
rect 619 103 627 108
rect 619 101 622 103
rect 624 101 627 103
rect 619 99 627 101
rect 629 110 637 117
rect 629 108 632 110
rect 634 108 637 110
rect 629 99 637 108
rect 639 120 644 126
rect 661 124 670 126
rect 661 122 663 124
rect 665 122 670 124
rect 639 118 646 120
rect 639 116 642 118
rect 644 116 646 118
rect 661 116 670 122
rect 639 114 646 116
rect 650 114 657 116
rect 639 99 644 114
rect 650 112 652 114
rect 654 112 657 114
rect 650 107 657 112
rect 650 105 652 107
rect 654 105 657 107
rect 650 103 657 105
rect 652 98 657 103
rect 659 105 670 116
rect 672 105 677 126
rect 679 119 684 126
rect 679 117 686 119
rect 701 117 707 119
rect 679 115 682 117
rect 684 115 686 117
rect 679 113 686 115
rect 679 105 684 113
rect 692 112 697 117
rect 690 110 697 112
rect 690 108 692 110
rect 694 108 697 110
rect 659 98 667 105
rect 690 103 697 108
rect 690 101 692 103
rect 694 101 697 103
rect 690 99 697 101
rect 699 115 707 117
rect 699 113 702 115
rect 704 113 707 115
rect 699 106 707 113
rect 709 117 717 119
rect 709 115 712 117
rect 714 115 717 117
rect 709 110 717 115
rect 709 108 712 110
rect 714 108 717 110
rect 709 106 717 108
rect 719 117 726 119
rect 719 115 722 117
rect 724 115 726 117
rect 719 106 726 115
rect 699 99 705 106
rect 741 105 746 126
rect 739 103 746 105
rect 739 101 741 103
rect 743 101 746 103
rect 739 99 746 101
rect 748 124 760 126
rect 748 122 751 124
rect 753 122 760 124
rect 748 117 760 122
rect 777 117 782 126
rect 748 115 751 117
rect 753 115 762 117
rect 748 99 762 115
rect 764 110 772 117
rect 764 108 767 110
rect 769 108 772 110
rect 764 103 772 108
rect 764 101 767 103
rect 769 101 772 103
rect 764 99 772 101
rect 774 110 782 117
rect 774 108 777 110
rect 779 108 782 110
rect 774 99 782 108
rect 784 120 789 126
rect 784 118 791 120
rect 784 116 787 118
rect 789 116 791 118
rect 806 117 812 119
rect 784 114 791 116
rect 784 99 789 114
rect 797 112 802 117
rect 795 110 802 112
rect 795 108 797 110
rect 799 108 802 110
rect 795 103 802 108
rect 795 101 797 103
rect 799 101 802 103
rect 795 99 802 101
rect 804 115 812 117
rect 804 113 807 115
rect 809 113 812 115
rect 804 106 812 113
rect 814 117 822 119
rect 814 115 817 117
rect 819 115 822 117
rect 814 110 822 115
rect 814 108 817 110
rect 819 108 822 110
rect 814 106 822 108
rect 824 117 831 119
rect 824 115 827 117
rect 829 115 831 117
rect 824 106 831 115
rect 804 99 810 106
rect 846 105 851 126
rect 844 103 851 105
rect 844 101 846 103
rect 848 101 851 103
rect 844 99 851 101
rect 853 124 865 126
rect 853 122 856 124
rect 858 122 865 124
rect 853 117 865 122
rect 882 117 887 126
rect 853 115 856 117
rect 858 115 867 117
rect 853 99 867 115
rect 869 110 877 117
rect 869 108 872 110
rect 874 108 877 110
rect 869 103 877 108
rect 869 101 872 103
rect 874 101 877 103
rect 869 99 877 101
rect 879 110 887 117
rect 879 108 882 110
rect 884 108 887 110
rect 879 99 887 108
rect 889 120 894 126
rect 911 124 920 126
rect 911 122 913 124
rect 915 122 920 124
rect 889 118 896 120
rect 889 116 892 118
rect 894 116 896 118
rect 911 116 920 122
rect 889 114 896 116
rect 900 114 907 116
rect 889 99 894 114
rect 900 112 902 114
rect 904 112 907 114
rect 900 107 907 112
rect 900 105 902 107
rect 904 105 907 107
rect 900 103 907 105
rect 902 98 907 103
rect 909 105 920 116
rect 922 105 927 126
rect 929 119 934 126
rect 929 117 936 119
rect 951 117 957 119
rect 929 115 932 117
rect 934 115 936 117
rect 929 113 936 115
rect 929 105 934 113
rect 942 112 947 117
rect 940 110 947 112
rect 940 108 942 110
rect 944 108 947 110
rect 909 98 917 105
rect 940 103 947 108
rect 940 101 942 103
rect 944 101 947 103
rect 940 99 947 101
rect 949 115 957 117
rect 949 113 952 115
rect 954 113 957 115
rect 949 106 957 113
rect 959 117 967 119
rect 959 115 962 117
rect 964 115 967 117
rect 959 110 967 115
rect 959 108 962 110
rect 964 108 967 110
rect 959 106 967 108
rect 969 117 976 119
rect 969 115 972 117
rect 974 115 976 117
rect 969 106 976 115
rect 949 99 955 106
rect 991 105 996 126
rect 989 103 996 105
rect 989 101 991 103
rect 993 101 996 103
rect 989 99 996 101
rect 998 124 1010 126
rect 998 122 1001 124
rect 1003 122 1010 124
rect 998 117 1010 122
rect 1027 117 1032 126
rect 998 115 1001 117
rect 1003 115 1012 117
rect 998 99 1012 115
rect 1014 110 1022 117
rect 1014 108 1017 110
rect 1019 108 1022 110
rect 1014 103 1022 108
rect 1014 101 1017 103
rect 1019 101 1022 103
rect 1014 99 1022 101
rect 1024 110 1032 117
rect 1024 108 1027 110
rect 1029 108 1032 110
rect 1024 99 1032 108
rect 1034 120 1039 126
rect 1034 118 1041 120
rect 1034 116 1037 118
rect 1039 116 1041 118
rect 1056 117 1062 119
rect 1034 114 1041 116
rect 1034 99 1039 114
rect 1047 112 1052 117
rect 1045 110 1052 112
rect 1045 108 1047 110
rect 1049 108 1052 110
rect 1045 103 1052 108
rect 1045 101 1047 103
rect 1049 101 1052 103
rect 1045 99 1052 101
rect 1054 115 1062 117
rect 1054 113 1057 115
rect 1059 113 1062 115
rect 1054 106 1062 113
rect 1064 117 1072 119
rect 1064 115 1067 117
rect 1069 115 1072 117
rect 1064 110 1072 115
rect 1064 108 1067 110
rect 1069 108 1072 110
rect 1064 106 1072 108
rect 1074 117 1081 119
rect 1074 115 1077 117
rect 1079 115 1081 117
rect 1074 106 1081 115
rect 1054 99 1060 106
rect 1096 105 1101 126
rect 1094 103 1101 105
rect 1094 101 1096 103
rect 1098 101 1101 103
rect 1094 99 1101 101
rect 1103 124 1115 126
rect 1103 122 1106 124
rect 1108 122 1115 124
rect 1103 117 1115 122
rect 1132 117 1137 126
rect 1103 115 1106 117
rect 1108 115 1117 117
rect 1103 99 1117 115
rect 1119 110 1127 117
rect 1119 108 1122 110
rect 1124 108 1127 110
rect 1119 103 1127 108
rect 1119 101 1122 103
rect 1124 101 1127 103
rect 1119 99 1127 101
rect 1129 110 1137 117
rect 1129 108 1132 110
rect 1134 108 1137 110
rect 1129 99 1137 108
rect 1139 120 1144 126
rect 1139 118 1146 120
rect 1139 116 1142 118
rect 1144 116 1146 118
rect 1139 114 1146 116
rect 1139 99 1144 114
rect 151 17 156 22
rect 149 15 156 17
rect 149 13 151 15
rect 153 13 156 15
rect 149 8 156 13
rect 149 6 151 8
rect 153 6 156 8
rect 149 4 156 6
rect 158 15 166 22
rect 189 19 196 21
rect 189 17 191 19
rect 193 17 196 19
rect 158 4 169 15
rect 160 -2 169 4
rect 160 -4 162 -2
rect 164 -4 169 -2
rect 160 -6 169 -4
rect 171 -6 176 15
rect 178 7 183 15
rect 189 12 196 17
rect 189 10 191 12
rect 193 10 196 12
rect 189 8 196 10
rect 178 5 185 7
rect 178 3 181 5
rect 183 3 185 5
rect 191 3 196 8
rect 198 14 204 21
rect 238 19 245 21
rect 238 17 240 19
rect 242 17 245 19
rect 238 15 245 17
rect 198 7 206 14
rect 198 5 201 7
rect 203 5 206 7
rect 198 3 206 5
rect 178 1 185 3
rect 178 -6 183 1
rect 200 1 206 3
rect 208 12 216 14
rect 208 10 211 12
rect 213 10 216 12
rect 208 5 216 10
rect 208 3 211 5
rect 213 3 216 5
rect 208 1 216 3
rect 218 5 225 14
rect 218 3 221 5
rect 223 3 225 5
rect 218 1 225 3
rect 240 -6 245 15
rect 247 5 261 21
rect 247 3 250 5
rect 252 3 261 5
rect 263 19 271 21
rect 263 17 266 19
rect 268 17 271 19
rect 263 12 271 17
rect 263 10 266 12
rect 268 10 271 12
rect 263 3 271 10
rect 273 12 281 21
rect 273 10 276 12
rect 278 10 281 12
rect 273 3 281 10
rect 247 -2 259 3
rect 247 -4 250 -2
rect 252 -4 259 -2
rect 247 -6 259 -4
rect 276 -6 281 3
rect 283 6 288 21
rect 294 19 301 21
rect 294 17 296 19
rect 298 17 301 19
rect 294 12 301 17
rect 294 10 296 12
rect 298 10 301 12
rect 294 8 301 10
rect 283 4 290 6
rect 283 2 286 4
rect 288 2 290 4
rect 296 3 301 8
rect 303 14 309 21
rect 343 19 350 21
rect 343 17 345 19
rect 347 17 350 19
rect 343 15 350 17
rect 303 7 311 14
rect 303 5 306 7
rect 308 5 311 7
rect 303 3 311 5
rect 283 0 290 2
rect 283 -6 288 0
rect 305 1 311 3
rect 313 12 321 14
rect 313 10 316 12
rect 318 10 321 12
rect 313 5 321 10
rect 313 3 316 5
rect 318 3 321 5
rect 313 1 321 3
rect 323 5 330 14
rect 323 3 326 5
rect 328 3 330 5
rect 323 1 330 3
rect 345 -6 350 15
rect 352 5 366 21
rect 352 3 355 5
rect 357 3 366 5
rect 368 19 376 21
rect 368 17 371 19
rect 373 17 376 19
rect 368 12 376 17
rect 368 10 371 12
rect 373 10 376 12
rect 368 3 376 10
rect 378 12 386 21
rect 378 10 381 12
rect 383 10 386 12
rect 378 3 386 10
rect 352 -2 364 3
rect 352 -4 355 -2
rect 357 -4 364 -2
rect 352 -6 364 -4
rect 381 -6 386 3
rect 388 6 393 21
rect 401 17 406 22
rect 399 15 406 17
rect 399 13 401 15
rect 403 13 406 15
rect 399 8 406 13
rect 399 6 401 8
rect 403 6 406 8
rect 388 4 395 6
rect 399 4 406 6
rect 408 15 416 22
rect 439 19 446 21
rect 439 17 441 19
rect 443 17 446 19
rect 408 4 419 15
rect 388 2 391 4
rect 393 2 395 4
rect 388 0 395 2
rect 388 -6 393 0
rect 410 -2 419 4
rect 410 -4 412 -2
rect 414 -4 419 -2
rect 410 -6 419 -4
rect 421 -6 426 15
rect 428 7 433 15
rect 439 12 446 17
rect 439 10 441 12
rect 443 10 446 12
rect 439 8 446 10
rect 428 5 435 7
rect 428 3 431 5
rect 433 3 435 5
rect 441 3 446 8
rect 448 14 454 21
rect 488 19 495 21
rect 488 17 490 19
rect 492 17 495 19
rect 488 15 495 17
rect 448 7 456 14
rect 448 5 451 7
rect 453 5 456 7
rect 448 3 456 5
rect 428 1 435 3
rect 428 -6 433 1
rect 450 1 456 3
rect 458 12 466 14
rect 458 10 461 12
rect 463 10 466 12
rect 458 5 466 10
rect 458 3 461 5
rect 463 3 466 5
rect 458 1 466 3
rect 468 5 475 14
rect 468 3 471 5
rect 473 3 475 5
rect 468 1 475 3
rect 490 -6 495 15
rect 497 5 511 21
rect 497 3 500 5
rect 502 3 511 5
rect 513 19 521 21
rect 513 17 516 19
rect 518 17 521 19
rect 513 12 521 17
rect 513 10 516 12
rect 518 10 521 12
rect 513 3 521 10
rect 523 12 531 21
rect 523 10 526 12
rect 528 10 531 12
rect 523 3 531 10
rect 497 -2 509 3
rect 497 -4 500 -2
rect 502 -4 509 -2
rect 497 -6 509 -4
rect 526 -6 531 3
rect 533 6 538 21
rect 544 19 551 21
rect 544 17 546 19
rect 548 17 551 19
rect 544 12 551 17
rect 544 10 546 12
rect 548 10 551 12
rect 544 8 551 10
rect 533 4 540 6
rect 533 2 536 4
rect 538 2 540 4
rect 546 3 551 8
rect 553 14 559 21
rect 593 19 600 21
rect 593 17 595 19
rect 597 17 600 19
rect 593 15 600 17
rect 553 7 561 14
rect 553 5 556 7
rect 558 5 561 7
rect 553 3 561 5
rect 533 0 540 2
rect 533 -6 538 0
rect 555 1 561 3
rect 563 12 571 14
rect 563 10 566 12
rect 568 10 571 12
rect 563 5 571 10
rect 563 3 566 5
rect 568 3 571 5
rect 563 1 571 3
rect 573 5 580 14
rect 573 3 576 5
rect 578 3 580 5
rect 573 1 580 3
rect 595 -6 600 15
rect 602 5 616 21
rect 602 3 605 5
rect 607 3 616 5
rect 618 19 626 21
rect 618 17 621 19
rect 623 17 626 19
rect 618 12 626 17
rect 618 10 621 12
rect 623 10 626 12
rect 618 3 626 10
rect 628 12 636 21
rect 628 10 631 12
rect 633 10 636 12
rect 628 3 636 10
rect 602 -2 614 3
rect 602 -4 605 -2
rect 607 -4 614 -2
rect 602 -6 614 -4
rect 631 -6 636 3
rect 638 6 643 21
rect 651 17 656 22
rect 649 15 656 17
rect 649 13 651 15
rect 653 13 656 15
rect 649 8 656 13
rect 649 6 651 8
rect 653 6 656 8
rect 638 4 645 6
rect 649 4 656 6
rect 658 15 666 22
rect 689 19 696 21
rect 689 17 691 19
rect 693 17 696 19
rect 658 4 669 15
rect 638 2 641 4
rect 643 2 645 4
rect 638 0 645 2
rect 638 -6 643 0
rect 660 -2 669 4
rect 660 -4 662 -2
rect 664 -4 669 -2
rect 660 -6 669 -4
rect 671 -6 676 15
rect 678 7 683 15
rect 689 12 696 17
rect 689 10 691 12
rect 693 10 696 12
rect 689 8 696 10
rect 678 5 685 7
rect 678 3 681 5
rect 683 3 685 5
rect 691 3 696 8
rect 698 14 704 21
rect 738 19 745 21
rect 738 17 740 19
rect 742 17 745 19
rect 738 15 745 17
rect 698 7 706 14
rect 698 5 701 7
rect 703 5 706 7
rect 698 3 706 5
rect 678 1 685 3
rect 678 -6 683 1
rect 700 1 706 3
rect 708 12 716 14
rect 708 10 711 12
rect 713 10 716 12
rect 708 5 716 10
rect 708 3 711 5
rect 713 3 716 5
rect 708 1 716 3
rect 718 5 725 14
rect 718 3 721 5
rect 723 3 725 5
rect 718 1 725 3
rect 740 -6 745 15
rect 747 5 761 21
rect 747 3 750 5
rect 752 3 761 5
rect 763 19 771 21
rect 763 17 766 19
rect 768 17 771 19
rect 763 12 771 17
rect 763 10 766 12
rect 768 10 771 12
rect 763 3 771 10
rect 773 12 781 21
rect 773 10 776 12
rect 778 10 781 12
rect 773 3 781 10
rect 747 -2 759 3
rect 747 -4 750 -2
rect 752 -4 759 -2
rect 747 -6 759 -4
rect 776 -6 781 3
rect 783 6 788 21
rect 794 19 801 21
rect 794 17 796 19
rect 798 17 801 19
rect 794 12 801 17
rect 794 10 796 12
rect 798 10 801 12
rect 794 8 801 10
rect 783 4 790 6
rect 783 2 786 4
rect 788 2 790 4
rect 796 3 801 8
rect 803 14 809 21
rect 843 19 850 21
rect 843 17 845 19
rect 847 17 850 19
rect 843 15 850 17
rect 803 7 811 14
rect 803 5 806 7
rect 808 5 811 7
rect 803 3 811 5
rect 783 0 790 2
rect 783 -6 788 0
rect 805 1 811 3
rect 813 12 821 14
rect 813 10 816 12
rect 818 10 821 12
rect 813 5 821 10
rect 813 3 816 5
rect 818 3 821 5
rect 813 1 821 3
rect 823 5 830 14
rect 823 3 826 5
rect 828 3 830 5
rect 823 1 830 3
rect 845 -6 850 15
rect 852 5 866 21
rect 852 3 855 5
rect 857 3 866 5
rect 868 19 876 21
rect 868 17 871 19
rect 873 17 876 19
rect 868 12 876 17
rect 868 10 871 12
rect 873 10 876 12
rect 868 3 876 10
rect 878 12 886 21
rect 878 10 881 12
rect 883 10 886 12
rect 878 3 886 10
rect 852 -2 864 3
rect 852 -4 855 -2
rect 857 -4 864 -2
rect 852 -6 864 -4
rect 881 -6 886 3
rect 888 6 893 21
rect 901 17 906 22
rect 899 15 906 17
rect 899 13 901 15
rect 903 13 906 15
rect 899 8 906 13
rect 899 6 901 8
rect 903 6 906 8
rect 888 4 895 6
rect 899 4 906 6
rect 908 15 916 22
rect 939 19 946 21
rect 939 17 941 19
rect 943 17 946 19
rect 908 4 919 15
rect 888 2 891 4
rect 893 2 895 4
rect 888 0 895 2
rect 888 -6 893 0
rect 910 -2 919 4
rect 910 -4 912 -2
rect 914 -4 919 -2
rect 910 -6 919 -4
rect 921 -6 926 15
rect 928 7 933 15
rect 939 12 946 17
rect 939 10 941 12
rect 943 10 946 12
rect 939 8 946 10
rect 928 5 935 7
rect 928 3 931 5
rect 933 3 935 5
rect 941 3 946 8
rect 948 14 954 21
rect 988 19 995 21
rect 988 17 990 19
rect 992 17 995 19
rect 988 15 995 17
rect 948 7 956 14
rect 948 5 951 7
rect 953 5 956 7
rect 948 3 956 5
rect 928 1 935 3
rect 928 -6 933 1
rect 950 1 956 3
rect 958 12 966 14
rect 958 10 961 12
rect 963 10 966 12
rect 958 5 966 10
rect 958 3 961 5
rect 963 3 966 5
rect 958 1 966 3
rect 968 5 975 14
rect 968 3 971 5
rect 973 3 975 5
rect 968 1 975 3
rect 990 -6 995 15
rect 997 5 1011 21
rect 997 3 1000 5
rect 1002 3 1011 5
rect 1013 19 1021 21
rect 1013 17 1016 19
rect 1018 17 1021 19
rect 1013 12 1021 17
rect 1013 10 1016 12
rect 1018 10 1021 12
rect 1013 3 1021 10
rect 1023 12 1031 21
rect 1023 10 1026 12
rect 1028 10 1031 12
rect 1023 3 1031 10
rect 997 -2 1009 3
rect 997 -4 1000 -2
rect 1002 -4 1009 -2
rect 997 -6 1009 -4
rect 1026 -6 1031 3
rect 1033 6 1038 21
rect 1044 19 1051 21
rect 1044 17 1046 19
rect 1048 17 1051 19
rect 1044 12 1051 17
rect 1044 10 1046 12
rect 1048 10 1051 12
rect 1044 8 1051 10
rect 1033 4 1040 6
rect 1033 2 1036 4
rect 1038 2 1040 4
rect 1046 3 1051 8
rect 1053 14 1059 21
rect 1093 19 1100 21
rect 1093 17 1095 19
rect 1097 17 1100 19
rect 1093 15 1100 17
rect 1053 7 1061 14
rect 1053 5 1056 7
rect 1058 5 1061 7
rect 1053 3 1061 5
rect 1033 0 1040 2
rect 1033 -6 1038 0
rect 1055 1 1061 3
rect 1063 12 1071 14
rect 1063 10 1066 12
rect 1068 10 1071 12
rect 1063 5 1071 10
rect 1063 3 1066 5
rect 1068 3 1071 5
rect 1063 1 1071 3
rect 1073 5 1080 14
rect 1073 3 1076 5
rect 1078 3 1080 5
rect 1073 1 1080 3
rect 1095 -6 1100 15
rect 1102 5 1116 21
rect 1102 3 1105 5
rect 1107 3 1116 5
rect 1118 19 1126 21
rect 1118 17 1121 19
rect 1123 17 1126 19
rect 1118 12 1126 17
rect 1118 10 1121 12
rect 1123 10 1126 12
rect 1118 3 1126 10
rect 1128 12 1136 21
rect 1128 10 1131 12
rect 1133 10 1136 12
rect 1128 3 1136 10
rect 1102 -2 1114 3
rect 1102 -4 1105 -2
rect 1107 -4 1114 -2
rect 1102 -6 1114 -4
rect 1131 -6 1136 3
rect 1138 6 1143 21
rect 1138 4 1145 6
rect 1138 2 1141 4
rect 1143 2 1145 4
rect 1138 0 1145 2
rect 1138 -6 1143 0
<< alu1 >>
rect 191 343 1029 348
rect 191 341 222 343
rect 224 341 232 343
rect 234 341 262 343
rect 264 341 272 343
rect 274 341 290 343
rect 292 341 343 343
rect 345 341 374 343
rect 376 341 384 343
rect 386 341 438 343
rect 440 341 448 343
rect 450 341 478 343
rect 480 341 488 343
rect 490 341 506 343
rect 508 341 559 343
rect 561 341 590 343
rect 592 341 600 343
rect 602 341 643 343
rect 645 341 653 343
rect 655 341 683 343
rect 685 341 693 343
rect 695 341 711 343
rect 713 341 764 343
rect 766 341 795 343
rect 797 341 805 343
rect 807 341 862 343
rect 864 341 872 343
rect 874 341 902 343
rect 904 341 912 343
rect 914 341 930 343
rect 932 341 983 343
rect 985 341 1014 343
rect 1016 341 1024 343
rect 1026 341 1029 343
rect 191 340 1029 341
rect 208 318 213 327
rect 225 331 237 335
rect 225 329 233 331
rect 235 329 237 331
rect 233 326 237 329
rect 208 317 222 318
rect 208 315 216 317
rect 218 315 219 317
rect 221 315 222 317
rect 208 314 222 315
rect 201 309 214 310
rect 201 307 206 309
rect 208 307 214 309
rect 201 306 214 307
rect 201 301 205 306
rect 233 324 234 326
rect 236 324 237 326
rect 233 309 237 324
rect 248 318 253 327
rect 265 331 277 335
rect 265 329 273 331
rect 275 329 277 331
rect 248 317 262 318
rect 248 315 256 317
rect 258 315 259 317
rect 261 315 262 317
rect 248 314 262 315
rect 201 299 202 301
rect 204 299 205 301
rect 201 297 205 299
rect 232 307 237 309
rect 232 305 233 307
rect 235 305 237 307
rect 232 300 237 305
rect 232 298 233 300
rect 235 298 237 300
rect 232 296 237 298
rect 241 309 254 310
rect 241 307 246 309
rect 248 307 254 309
rect 241 306 254 307
rect 241 302 245 306
rect 273 309 277 329
rect 241 300 242 302
rect 244 300 245 302
rect 241 297 245 300
rect 272 307 277 309
rect 272 305 273 307
rect 275 305 277 307
rect 272 303 277 305
rect 272 301 273 303
rect 275 301 277 303
rect 272 300 277 301
rect 272 298 273 300
rect 275 298 277 300
rect 272 296 277 298
rect 288 333 312 334
rect 288 331 308 333
rect 310 331 312 333
rect 288 330 312 331
rect 288 302 292 330
rect 327 326 340 327
rect 327 324 335 326
rect 337 324 340 326
rect 327 322 340 324
rect 327 320 328 322
rect 330 321 340 322
rect 330 320 332 321
rect 288 300 304 302
rect 288 298 300 300
rect 302 298 304 300
rect 288 297 304 298
rect 327 313 332 320
rect 360 326 365 327
rect 360 324 362 326
rect 364 324 365 326
rect 360 318 365 324
rect 377 331 389 335
rect 377 329 385 331
rect 387 329 389 331
rect 360 317 374 318
rect 360 315 368 317
rect 370 315 374 317
rect 360 314 374 315
rect 343 310 348 311
rect 343 309 349 310
rect 353 309 366 310
rect 343 307 344 309
rect 346 307 358 309
rect 360 307 366 309
rect 343 306 366 307
rect 343 304 357 306
rect 343 295 348 304
rect 353 303 357 304
rect 385 314 389 329
rect 424 318 429 327
rect 441 331 453 335
rect 441 329 449 331
rect 451 329 453 331
rect 449 326 453 329
rect 424 317 438 318
rect 424 315 432 317
rect 434 315 435 317
rect 437 315 438 317
rect 424 314 438 315
rect 385 312 386 314
rect 388 312 389 314
rect 385 309 389 312
rect 353 301 354 303
rect 356 301 357 303
rect 353 297 357 301
rect 384 307 389 309
rect 384 305 385 307
rect 387 305 389 307
rect 384 300 389 305
rect 336 289 348 295
rect 384 298 385 300
rect 387 298 389 300
rect 384 296 389 298
rect 417 309 430 310
rect 417 307 422 309
rect 424 307 430 309
rect 417 306 430 307
rect 417 301 421 306
rect 449 324 450 326
rect 452 324 453 326
rect 449 309 453 324
rect 464 318 469 327
rect 481 331 493 335
rect 481 329 489 331
rect 491 329 493 331
rect 464 317 478 318
rect 464 315 472 317
rect 474 315 475 317
rect 477 315 478 317
rect 464 314 478 315
rect 417 299 418 301
rect 420 299 421 301
rect 417 297 421 299
rect 448 307 453 309
rect 448 305 449 307
rect 451 305 453 307
rect 448 300 453 305
rect 448 298 449 300
rect 451 298 453 300
rect 448 296 453 298
rect 457 309 470 310
rect 457 307 462 309
rect 464 307 470 309
rect 457 306 470 307
rect 457 302 461 306
rect 489 309 493 329
rect 457 300 458 302
rect 460 300 461 302
rect 457 297 461 300
rect 488 307 493 309
rect 488 305 489 307
rect 491 305 493 307
rect 488 303 493 305
rect 488 301 489 303
rect 491 301 493 303
rect 488 300 493 301
rect 488 298 489 300
rect 491 298 493 300
rect 488 296 493 298
rect 504 333 528 334
rect 504 331 524 333
rect 526 331 528 333
rect 504 330 528 331
rect 504 302 508 330
rect 543 326 556 327
rect 543 324 551 326
rect 553 324 556 326
rect 543 322 556 324
rect 543 320 544 322
rect 546 321 556 322
rect 546 320 548 321
rect 504 300 520 302
rect 504 298 516 300
rect 518 298 520 300
rect 504 297 520 298
rect 543 313 548 320
rect 576 326 581 327
rect 576 324 578 326
rect 580 324 581 326
rect 576 318 581 324
rect 593 331 605 335
rect 593 329 601 331
rect 603 329 605 331
rect 576 317 590 318
rect 576 315 584 317
rect 586 315 590 317
rect 576 314 590 315
rect 559 310 564 311
rect 559 309 565 310
rect 569 309 582 310
rect 559 307 560 309
rect 562 307 574 309
rect 576 307 582 309
rect 559 306 582 307
rect 559 304 573 306
rect 559 295 564 304
rect 569 303 573 304
rect 601 314 605 329
rect 629 318 634 327
rect 646 331 658 335
rect 646 329 654 331
rect 656 329 658 331
rect 654 326 658 329
rect 629 317 643 318
rect 629 315 637 317
rect 639 315 640 317
rect 642 315 643 317
rect 629 314 643 315
rect 601 312 602 314
rect 604 312 605 314
rect 601 309 605 312
rect 569 301 570 303
rect 572 301 573 303
rect 569 297 573 301
rect 600 307 605 309
rect 600 305 601 307
rect 603 305 605 307
rect 600 300 605 305
rect 552 289 564 295
rect 600 298 601 300
rect 603 298 605 300
rect 600 296 605 298
rect 622 309 635 310
rect 622 307 627 309
rect 629 307 635 309
rect 622 306 635 307
rect 622 301 626 306
rect 654 324 655 326
rect 657 324 658 326
rect 654 309 658 324
rect 669 318 674 327
rect 686 331 698 335
rect 686 329 694 331
rect 696 329 698 331
rect 669 317 683 318
rect 669 315 677 317
rect 679 315 680 317
rect 682 315 683 317
rect 669 314 683 315
rect 622 299 623 301
rect 625 299 626 301
rect 622 297 626 299
rect 653 307 658 309
rect 653 305 654 307
rect 656 305 658 307
rect 653 300 658 305
rect 653 298 654 300
rect 656 298 658 300
rect 653 296 658 298
rect 662 309 675 310
rect 662 307 667 309
rect 669 307 675 309
rect 662 306 675 307
rect 662 302 666 306
rect 694 309 698 329
rect 662 300 663 302
rect 665 300 666 302
rect 662 297 666 300
rect 693 307 698 309
rect 693 305 694 307
rect 696 305 698 307
rect 693 303 698 305
rect 693 301 694 303
rect 696 301 698 303
rect 693 300 698 301
rect 693 298 694 300
rect 696 298 698 300
rect 693 296 698 298
rect 709 333 733 334
rect 709 331 729 333
rect 731 331 733 333
rect 709 330 733 331
rect 709 302 713 330
rect 748 326 761 327
rect 748 324 756 326
rect 758 324 761 326
rect 748 322 761 324
rect 748 320 749 322
rect 751 321 761 322
rect 751 320 753 321
rect 709 300 725 302
rect 709 298 721 300
rect 723 298 725 300
rect 709 297 725 298
rect 748 313 753 320
rect 781 326 786 327
rect 781 324 783 326
rect 785 324 786 326
rect 781 318 786 324
rect 798 331 810 335
rect 798 329 806 331
rect 808 329 810 331
rect 781 317 795 318
rect 781 315 789 317
rect 791 315 795 317
rect 781 314 795 315
rect 764 310 769 311
rect 764 309 770 310
rect 774 309 787 310
rect 764 307 765 309
rect 767 307 779 309
rect 781 307 787 309
rect 764 306 787 307
rect 764 304 778 306
rect 764 295 769 304
rect 774 303 778 304
rect 806 314 810 329
rect 848 318 853 327
rect 865 331 877 335
rect 865 329 873 331
rect 875 329 877 331
rect 873 326 877 329
rect 848 317 862 318
rect 848 315 856 317
rect 858 315 859 317
rect 861 315 862 317
rect 848 314 862 315
rect 806 312 807 314
rect 809 312 810 314
rect 806 309 810 312
rect 774 301 775 303
rect 777 301 778 303
rect 774 297 778 301
rect 805 307 810 309
rect 805 305 806 307
rect 808 305 810 307
rect 805 300 810 305
rect 757 289 769 295
rect 805 298 806 300
rect 808 298 810 300
rect 805 296 810 298
rect 841 309 854 310
rect 841 307 846 309
rect 848 307 854 309
rect 841 306 854 307
rect 841 301 845 306
rect 873 324 874 326
rect 876 324 877 326
rect 873 309 877 324
rect 888 318 893 327
rect 905 331 917 335
rect 905 329 913 331
rect 915 329 917 331
rect 888 317 902 318
rect 888 315 896 317
rect 898 315 899 317
rect 901 315 902 317
rect 888 314 902 315
rect 841 299 842 301
rect 844 299 845 301
rect 841 297 845 299
rect 872 307 877 309
rect 872 305 873 307
rect 875 305 877 307
rect 872 300 877 305
rect 872 298 873 300
rect 875 298 877 300
rect 872 296 877 298
rect 881 309 894 310
rect 881 307 886 309
rect 888 307 894 309
rect 881 306 894 307
rect 881 302 885 306
rect 913 309 917 329
rect 881 300 882 302
rect 884 300 885 302
rect 881 297 885 300
rect 912 307 917 309
rect 912 305 913 307
rect 915 305 917 307
rect 912 303 917 305
rect 912 301 913 303
rect 915 301 917 303
rect 912 300 917 301
rect 912 298 913 300
rect 915 298 917 300
rect 912 296 917 298
rect 928 333 952 334
rect 928 331 948 333
rect 950 331 952 333
rect 928 330 952 331
rect 928 302 932 330
rect 967 326 980 327
rect 967 324 975 326
rect 977 324 980 326
rect 967 322 980 324
rect 967 320 968 322
rect 970 321 980 322
rect 970 320 972 321
rect 928 300 944 302
rect 928 298 940 300
rect 942 298 944 300
rect 928 297 944 298
rect 967 313 972 320
rect 1000 326 1005 327
rect 1000 324 1002 326
rect 1004 324 1005 326
rect 1000 318 1005 324
rect 1017 331 1029 335
rect 1017 329 1025 331
rect 1027 329 1029 331
rect 1000 317 1014 318
rect 1000 315 1008 317
rect 1010 315 1014 317
rect 1000 314 1014 315
rect 983 310 988 311
rect 983 309 989 310
rect 993 309 1006 310
rect 983 307 984 309
rect 986 307 998 309
rect 1000 307 1006 309
rect 983 306 1006 307
rect 983 304 997 306
rect 983 295 988 304
rect 993 303 997 304
rect 1025 314 1029 329
rect 1025 312 1026 314
rect 1028 312 1029 314
rect 1025 309 1029 312
rect 993 301 994 303
rect 996 301 997 303
rect 993 297 997 301
rect 1024 307 1029 309
rect 1024 305 1025 307
rect 1027 305 1029 307
rect 1024 300 1029 305
rect 976 289 988 295
rect 1024 298 1025 300
rect 1027 298 1029 300
rect 1024 296 1029 298
rect 200 283 389 284
rect 200 281 232 283
rect 234 281 272 283
rect 274 281 310 283
rect 312 281 384 283
rect 386 281 389 283
rect 200 271 389 281
rect 200 269 204 271
rect 206 269 272 271
rect 274 269 284 271
rect 286 269 358 271
rect 360 269 389 271
rect 200 268 389 269
rect 416 283 810 284
rect 416 281 448 283
rect 450 281 488 283
rect 490 281 526 283
rect 528 281 600 283
rect 602 281 653 283
rect 655 281 693 283
rect 695 281 731 283
rect 733 281 805 283
rect 807 281 810 283
rect 416 271 810 281
rect 416 269 420 271
rect 422 269 488 271
rect 490 269 500 271
rect 502 269 574 271
rect 576 269 625 271
rect 627 269 693 271
rect 695 269 705 271
rect 707 269 779 271
rect 781 269 810 271
rect 416 268 810 269
rect 840 283 1029 284
rect 840 281 872 283
rect 874 281 912 283
rect 914 281 950 283
rect 952 281 1024 283
rect 1026 281 1029 283
rect 840 271 1029 281
rect 840 269 844 271
rect 846 269 912 271
rect 914 269 924 271
rect 926 269 998 271
rect 1000 269 1029 271
rect 840 268 1029 269
rect 1041 271 1150 276
rect 1041 269 1048 271
rect 1050 269 1122 271
rect 1124 269 1150 271
rect 1041 268 1150 269
rect 201 254 206 256
rect 201 252 203 254
rect 205 252 206 254
rect 201 247 206 252
rect 201 245 203 247
rect 205 245 206 247
rect 201 243 206 245
rect 233 254 237 255
rect 233 252 234 254
rect 236 252 237 254
rect 201 223 205 243
rect 233 246 237 252
rect 224 245 237 246
rect 224 243 230 245
rect 232 243 237 245
rect 224 242 237 243
rect 241 246 245 255
rect 272 254 277 256
rect 241 245 254 246
rect 241 243 242 245
rect 244 243 246 245
rect 248 243 254 245
rect 241 242 254 243
rect 216 237 230 238
rect 216 235 217 237
rect 219 235 220 237
rect 222 235 230 237
rect 216 234 230 235
rect 201 221 203 223
rect 205 221 213 223
rect 201 217 213 221
rect 225 225 230 234
rect 248 237 262 238
rect 248 235 256 237
rect 258 235 259 237
rect 261 235 262 237
rect 248 234 262 235
rect 272 252 273 254
rect 275 252 277 254
rect 272 247 277 252
rect 272 245 273 247
rect 275 245 277 247
rect 272 243 277 245
rect 248 225 253 234
rect 273 228 277 243
rect 273 226 274 228
rect 276 226 277 228
rect 273 223 277 226
rect 265 221 273 223
rect 275 221 277 223
rect 265 217 277 221
rect 281 254 286 256
rect 281 252 283 254
rect 285 252 286 254
rect 322 261 334 263
rect 322 259 330 261
rect 332 259 334 261
rect 322 257 334 259
rect 281 247 286 252
rect 281 245 283 247
rect 285 245 286 247
rect 281 243 286 245
rect 281 223 285 243
rect 313 248 317 255
rect 322 248 327 257
rect 313 246 327 248
rect 304 245 327 246
rect 304 243 310 245
rect 312 243 324 245
rect 326 243 327 245
rect 304 242 317 243
rect 321 242 327 243
rect 322 241 327 242
rect 296 237 310 238
rect 296 235 300 237
rect 302 235 310 237
rect 296 234 310 235
rect 281 221 283 223
rect 285 221 293 223
rect 281 217 293 221
rect 305 228 310 234
rect 305 226 306 228
rect 308 226 310 228
rect 305 225 310 226
rect 338 232 343 239
rect 366 254 382 255
rect 366 252 368 254
rect 370 252 382 254
rect 366 250 382 252
rect 338 231 340 232
rect 330 230 340 231
rect 342 230 343 232
rect 330 228 343 230
rect 330 226 333 228
rect 335 226 343 228
rect 330 225 343 226
rect 378 222 382 250
rect 358 221 382 222
rect 358 219 360 221
rect 362 219 382 221
rect 358 218 382 219
rect 417 254 422 256
rect 417 252 419 254
rect 421 252 422 254
rect 417 247 422 252
rect 417 245 419 247
rect 421 245 422 247
rect 417 243 422 245
rect 449 254 453 255
rect 449 252 450 254
rect 452 252 453 254
rect 417 223 421 243
rect 449 246 453 252
rect 440 245 453 246
rect 440 243 446 245
rect 448 243 453 245
rect 440 242 453 243
rect 457 246 461 255
rect 488 254 493 256
rect 457 245 470 246
rect 457 243 458 245
rect 460 243 462 245
rect 464 243 470 245
rect 457 242 470 243
rect 432 237 446 238
rect 432 235 433 237
rect 435 235 436 237
rect 438 235 446 237
rect 432 234 446 235
rect 417 221 419 223
rect 421 221 429 223
rect 417 217 429 221
rect 441 225 446 234
rect 464 237 478 238
rect 464 235 472 237
rect 474 235 475 237
rect 477 235 478 237
rect 464 234 478 235
rect 488 252 489 254
rect 491 252 493 254
rect 488 247 493 252
rect 488 245 489 247
rect 491 245 493 247
rect 488 243 493 245
rect 464 225 469 234
rect 489 228 493 243
rect 489 226 490 228
rect 492 226 493 228
rect 489 223 493 226
rect 481 221 489 223
rect 491 221 493 223
rect 481 217 493 221
rect 497 254 502 256
rect 497 252 499 254
rect 501 252 502 254
rect 538 261 550 263
rect 538 259 546 261
rect 548 259 550 261
rect 538 257 550 259
rect 497 247 502 252
rect 497 245 499 247
rect 501 245 502 247
rect 497 243 502 245
rect 497 223 501 243
rect 529 248 533 255
rect 538 248 543 257
rect 529 246 543 248
rect 520 245 543 246
rect 520 243 526 245
rect 528 243 540 245
rect 542 243 543 245
rect 520 242 533 243
rect 537 242 543 243
rect 538 241 543 242
rect 512 237 526 238
rect 512 235 516 237
rect 518 235 526 237
rect 512 234 526 235
rect 497 221 499 223
rect 501 221 509 223
rect 497 217 509 221
rect 521 228 526 234
rect 521 226 522 228
rect 524 226 526 228
rect 521 225 526 226
rect 554 232 559 239
rect 582 254 598 255
rect 582 252 584 254
rect 586 252 598 254
rect 582 250 598 252
rect 554 231 556 232
rect 546 230 556 231
rect 558 230 559 232
rect 546 228 559 230
rect 546 226 549 228
rect 551 226 559 228
rect 546 225 559 226
rect 594 222 598 250
rect 574 221 598 222
rect 574 219 576 221
rect 578 219 598 221
rect 574 218 598 219
rect 622 254 627 256
rect 622 252 624 254
rect 626 252 627 254
rect 622 247 627 252
rect 622 245 624 247
rect 626 245 627 247
rect 622 243 627 245
rect 654 254 658 255
rect 654 252 655 254
rect 657 252 658 254
rect 622 223 626 243
rect 654 246 658 252
rect 645 245 658 246
rect 645 243 651 245
rect 653 243 658 245
rect 645 242 658 243
rect 662 246 666 255
rect 693 254 698 256
rect 662 245 675 246
rect 662 243 663 245
rect 665 243 667 245
rect 669 243 675 245
rect 662 242 675 243
rect 637 237 651 238
rect 637 235 638 237
rect 640 235 641 237
rect 643 235 651 237
rect 637 234 651 235
rect 622 221 624 223
rect 626 221 634 223
rect 622 217 634 221
rect 646 225 651 234
rect 669 237 683 238
rect 669 235 677 237
rect 679 235 680 237
rect 682 235 683 237
rect 669 234 683 235
rect 693 252 694 254
rect 696 252 698 254
rect 693 247 698 252
rect 693 245 694 247
rect 696 245 698 247
rect 693 243 698 245
rect 669 225 674 234
rect 694 228 698 243
rect 694 226 695 228
rect 697 226 698 228
rect 694 223 698 226
rect 686 221 694 223
rect 696 221 698 223
rect 686 217 698 221
rect 702 254 707 256
rect 702 252 704 254
rect 706 252 707 254
rect 743 261 755 263
rect 743 259 751 261
rect 753 259 755 261
rect 743 257 755 259
rect 702 247 707 252
rect 702 245 704 247
rect 706 245 707 247
rect 702 243 707 245
rect 702 223 706 243
rect 734 248 738 255
rect 743 248 748 257
rect 734 246 748 248
rect 725 245 748 246
rect 725 243 731 245
rect 733 243 745 245
rect 747 243 748 245
rect 725 242 738 243
rect 742 242 748 243
rect 743 241 748 242
rect 717 237 731 238
rect 717 235 721 237
rect 723 235 731 237
rect 717 234 731 235
rect 702 221 704 223
rect 706 221 714 223
rect 702 217 714 221
rect 726 228 731 234
rect 726 226 727 228
rect 729 226 731 228
rect 726 225 731 226
rect 759 232 764 239
rect 787 254 803 255
rect 787 252 789 254
rect 791 252 803 254
rect 787 250 803 252
rect 759 231 761 232
rect 751 230 761 231
rect 763 230 764 232
rect 751 228 764 230
rect 751 226 754 228
rect 756 226 764 228
rect 751 225 764 226
rect 799 222 803 250
rect 779 221 803 222
rect 779 219 781 221
rect 783 219 803 221
rect 779 218 803 219
rect 841 254 846 256
rect 841 252 843 254
rect 845 252 846 254
rect 841 247 846 252
rect 841 245 843 247
rect 845 245 846 247
rect 841 243 846 245
rect 873 254 877 255
rect 873 252 874 254
rect 876 252 877 254
rect 841 223 845 243
rect 873 246 877 252
rect 864 245 877 246
rect 864 243 870 245
rect 872 243 877 245
rect 864 242 877 243
rect 881 246 885 255
rect 912 254 917 256
rect 881 245 894 246
rect 881 243 882 245
rect 884 243 886 245
rect 888 243 894 245
rect 881 242 894 243
rect 856 237 870 238
rect 856 235 857 237
rect 859 235 860 237
rect 862 235 870 237
rect 856 234 870 235
rect 841 221 843 223
rect 845 221 853 223
rect 841 217 853 221
rect 865 225 870 234
rect 888 237 902 238
rect 888 235 896 237
rect 898 235 899 237
rect 901 235 902 237
rect 888 234 902 235
rect 912 252 913 254
rect 915 252 917 254
rect 912 247 917 252
rect 912 245 913 247
rect 915 245 917 247
rect 912 243 917 245
rect 888 225 893 234
rect 913 228 917 243
rect 913 226 914 228
rect 916 226 917 228
rect 913 223 917 226
rect 905 221 913 223
rect 915 221 917 223
rect 905 217 917 221
rect 921 254 926 256
rect 921 252 923 254
rect 925 252 926 254
rect 962 261 974 263
rect 962 259 970 261
rect 972 259 974 261
rect 962 257 974 259
rect 921 247 926 252
rect 921 245 923 247
rect 925 245 926 247
rect 921 243 926 245
rect 921 223 925 243
rect 953 248 957 255
rect 962 248 967 257
rect 953 246 967 248
rect 944 245 967 246
rect 944 243 950 245
rect 952 243 964 245
rect 966 243 967 245
rect 944 242 957 243
rect 961 242 967 243
rect 962 241 967 242
rect 936 237 950 238
rect 936 235 940 237
rect 942 235 950 237
rect 936 234 950 235
rect 921 221 923 223
rect 925 221 933 223
rect 921 217 933 221
rect 945 228 950 234
rect 945 226 946 228
rect 948 226 950 228
rect 945 225 950 226
rect 978 232 983 239
rect 1006 254 1022 255
rect 1006 252 1008 254
rect 1010 252 1022 254
rect 1006 250 1022 252
rect 978 231 980 232
rect 970 230 980 231
rect 982 230 983 232
rect 970 228 983 230
rect 970 226 973 228
rect 975 226 983 228
rect 970 225 983 226
rect 1018 222 1022 250
rect 998 221 1022 222
rect 998 219 1000 221
rect 1002 219 1022 221
rect 998 218 1022 219
rect 1045 254 1050 256
rect 1045 252 1047 254
rect 1049 252 1050 254
rect 1086 257 1098 263
rect 1045 247 1050 252
rect 1045 245 1047 247
rect 1049 245 1050 247
rect 1045 243 1050 245
rect 1045 223 1049 243
rect 1077 248 1081 255
rect 1086 248 1091 257
rect 1077 246 1091 248
rect 1068 245 1091 246
rect 1068 243 1074 245
rect 1076 243 1088 245
rect 1090 243 1091 245
rect 1068 242 1081 243
rect 1085 242 1091 243
rect 1086 241 1091 242
rect 1060 237 1074 238
rect 1060 235 1064 237
rect 1066 235 1074 237
rect 1060 234 1074 235
rect 1045 221 1047 223
rect 1049 221 1057 223
rect 1045 217 1057 221
rect 1069 228 1074 234
rect 1069 226 1070 228
rect 1072 226 1074 228
rect 1069 225 1074 226
rect 1102 232 1107 239
rect 1130 254 1146 255
rect 1130 252 1132 254
rect 1134 252 1146 254
rect 1130 250 1146 252
rect 1102 231 1104 232
rect 1094 230 1104 231
rect 1106 230 1107 232
rect 1094 228 1107 230
rect 1094 226 1097 228
rect 1099 226 1107 228
rect 1094 225 1107 226
rect 1142 222 1146 250
rect 1122 221 1146 222
rect 1122 219 1124 221
rect 1126 219 1146 221
rect 1122 218 1146 219
rect 191 211 1026 212
rect 191 209 204 211
rect 206 209 214 211
rect 216 209 262 211
rect 264 209 272 211
rect 274 209 284 211
rect 286 209 294 211
rect 296 209 325 211
rect 327 209 378 211
rect 380 209 420 211
rect 422 209 430 211
rect 432 209 478 211
rect 480 209 488 211
rect 490 209 500 211
rect 502 209 510 211
rect 512 209 541 211
rect 543 209 594 211
rect 596 209 625 211
rect 627 209 635 211
rect 637 209 683 211
rect 685 209 693 211
rect 695 209 705 211
rect 707 209 715 211
rect 717 209 746 211
rect 748 209 799 211
rect 801 209 844 211
rect 846 209 854 211
rect 856 209 902 211
rect 904 209 912 211
rect 914 209 924 211
rect 926 209 934 211
rect 936 209 965 211
rect 967 209 1018 211
rect 1020 209 1026 211
rect 191 204 1026 209
rect 1041 211 1150 212
rect 1041 209 1048 211
rect 1050 209 1058 211
rect 1060 209 1089 211
rect 1091 209 1142 211
rect 1144 209 1150 211
rect 1041 204 1150 209
rect 147 199 1151 204
rect 147 197 154 199
rect 156 197 194 199
rect 196 197 204 199
rect 206 197 235 199
rect 237 197 288 199
rect 290 197 299 199
rect 301 197 309 199
rect 311 197 340 199
rect 342 197 393 199
rect 395 197 404 199
rect 406 197 444 199
rect 446 197 454 199
rect 456 197 485 199
rect 487 197 538 199
rect 540 197 549 199
rect 551 197 559 199
rect 561 197 590 199
rect 592 197 643 199
rect 645 197 654 199
rect 656 197 694 199
rect 696 197 704 199
rect 706 197 735 199
rect 737 197 788 199
rect 790 197 799 199
rect 801 197 809 199
rect 811 197 840 199
rect 842 197 893 199
rect 895 197 904 199
rect 906 197 944 199
rect 946 197 954 199
rect 956 197 985 199
rect 987 197 1038 199
rect 1040 197 1049 199
rect 1051 197 1059 199
rect 1061 197 1090 199
rect 1092 197 1143 199
rect 1145 197 1151 199
rect 147 196 1151 197
rect 191 187 203 191
rect 191 185 193 187
rect 195 185 203 187
rect 268 189 292 190
rect 151 182 156 184
rect 151 180 153 182
rect 155 180 156 182
rect 151 178 156 180
rect 151 159 155 178
rect 183 174 187 183
rect 191 174 195 185
rect 268 187 270 189
rect 272 187 292 189
rect 268 186 292 187
rect 151 157 153 159
rect 151 152 155 157
rect 151 150 153 152
rect 166 173 195 174
rect 166 171 170 173
rect 172 171 195 173
rect 166 170 195 171
rect 166 164 180 166
rect 182 164 187 166
rect 166 162 187 164
rect 183 156 187 162
rect 183 154 184 156
rect 186 154 187 156
rect 183 153 187 154
rect 191 165 195 170
rect 215 182 220 183
rect 215 180 216 182
rect 218 180 220 182
rect 215 174 220 180
rect 191 163 196 165
rect 191 161 193 163
rect 195 161 196 163
rect 191 156 196 161
rect 191 154 193 156
rect 195 154 196 156
rect 206 173 220 174
rect 206 171 210 173
rect 212 171 220 173
rect 206 170 220 171
rect 240 182 253 183
rect 240 180 243 182
rect 245 180 253 182
rect 240 178 253 180
rect 288 182 292 186
rect 240 177 250 178
rect 248 176 250 177
rect 252 176 253 178
rect 232 166 237 167
rect 214 165 227 166
rect 231 165 237 166
rect 214 163 220 165
rect 222 163 234 165
rect 236 163 237 165
rect 214 162 237 163
rect 223 160 237 162
rect 248 169 253 176
rect 288 180 289 182
rect 291 180 292 182
rect 191 152 196 154
rect 151 146 164 150
rect 151 145 155 146
rect 223 153 227 160
rect 232 151 237 160
rect 232 145 244 151
rect 288 158 292 180
rect 276 156 292 158
rect 276 154 278 156
rect 280 154 292 156
rect 276 153 292 154
rect 296 187 308 191
rect 296 185 298 187
rect 300 185 308 187
rect 373 189 397 190
rect 296 165 300 185
rect 373 187 375 189
rect 377 187 397 189
rect 373 186 397 187
rect 320 182 325 183
rect 320 180 321 182
rect 323 180 325 182
rect 320 174 325 180
rect 296 163 301 165
rect 296 161 298 163
rect 300 161 301 163
rect 296 156 301 161
rect 296 154 298 156
rect 300 154 301 156
rect 311 173 325 174
rect 311 171 315 173
rect 317 171 325 173
rect 311 170 325 171
rect 345 182 358 183
rect 345 180 348 182
rect 350 180 358 182
rect 345 178 358 180
rect 345 177 355 178
rect 353 176 355 177
rect 357 176 358 178
rect 337 166 342 167
rect 319 165 332 166
rect 336 165 342 166
rect 319 163 325 165
rect 327 164 339 165
rect 327 163 331 164
rect 319 162 331 163
rect 333 163 339 164
rect 341 163 342 165
rect 333 162 342 163
rect 328 160 342 162
rect 353 169 358 176
rect 296 152 301 154
rect 328 153 332 160
rect 337 151 342 160
rect 337 145 349 151
rect 393 158 397 186
rect 441 187 453 191
rect 441 185 443 187
rect 445 185 453 187
rect 518 189 542 190
rect 381 156 397 158
rect 381 154 383 156
rect 385 154 397 156
rect 381 153 397 154
rect 401 182 406 184
rect 401 180 403 182
rect 405 180 406 182
rect 401 178 406 180
rect 401 164 405 178
rect 401 162 402 164
rect 404 162 405 164
rect 401 159 405 162
rect 433 174 437 183
rect 441 174 445 185
rect 518 187 520 189
rect 522 187 542 189
rect 518 186 542 187
rect 401 157 403 159
rect 401 152 405 157
rect 401 150 403 152
rect 416 173 445 174
rect 416 171 420 173
rect 422 171 445 173
rect 416 170 445 171
rect 416 164 430 166
rect 432 164 437 166
rect 416 162 437 164
rect 433 156 437 162
rect 433 154 434 156
rect 436 154 437 156
rect 433 153 437 154
rect 441 165 445 170
rect 465 182 470 183
rect 465 180 466 182
rect 468 180 470 182
rect 465 174 470 180
rect 441 163 446 165
rect 441 161 443 163
rect 445 161 446 163
rect 441 156 446 161
rect 441 154 443 156
rect 445 154 446 156
rect 456 173 470 174
rect 456 171 460 173
rect 462 171 470 173
rect 456 170 470 171
rect 490 182 503 183
rect 490 180 493 182
rect 495 180 503 182
rect 490 178 503 180
rect 538 182 542 186
rect 490 177 500 178
rect 498 176 500 177
rect 502 176 503 178
rect 482 166 487 167
rect 464 165 477 166
rect 481 165 487 166
rect 464 163 470 165
rect 472 163 484 165
rect 486 163 487 165
rect 464 162 487 163
rect 473 160 487 162
rect 498 169 503 176
rect 538 180 539 182
rect 541 180 542 182
rect 441 152 446 154
rect 401 146 414 150
rect 401 145 405 146
rect 473 153 477 160
rect 482 151 487 160
rect 482 145 494 151
rect 538 158 542 180
rect 526 156 542 158
rect 526 154 528 156
rect 530 154 542 156
rect 526 153 542 154
rect 546 187 558 191
rect 546 185 548 187
rect 550 185 558 187
rect 623 189 647 190
rect 546 165 550 185
rect 623 187 625 189
rect 627 187 647 189
rect 623 186 647 187
rect 570 182 575 183
rect 570 180 571 182
rect 573 180 575 182
rect 570 174 575 180
rect 546 163 551 165
rect 546 161 548 163
rect 550 161 551 163
rect 546 156 551 161
rect 546 154 548 156
rect 550 154 551 156
rect 561 173 575 174
rect 561 171 565 173
rect 567 171 575 173
rect 561 170 575 171
rect 595 182 608 183
rect 595 180 598 182
rect 600 180 608 182
rect 595 178 608 180
rect 595 177 605 178
rect 603 176 605 177
rect 607 176 608 178
rect 587 166 592 167
rect 569 165 582 166
rect 586 165 592 166
rect 569 163 575 165
rect 577 164 589 165
rect 577 163 583 164
rect 569 162 583 163
rect 585 163 589 164
rect 591 163 592 165
rect 585 162 592 163
rect 578 160 592 162
rect 603 169 608 176
rect 546 152 551 154
rect 578 153 582 160
rect 587 151 592 160
rect 587 145 599 151
rect 643 158 647 186
rect 691 187 703 191
rect 691 185 693 187
rect 695 185 703 187
rect 768 189 792 190
rect 631 156 647 158
rect 631 154 633 156
rect 635 154 647 156
rect 631 153 647 154
rect 651 182 656 184
rect 651 180 653 182
rect 655 180 656 182
rect 651 178 656 180
rect 651 164 655 178
rect 651 162 652 164
rect 654 162 655 164
rect 651 159 655 162
rect 683 174 687 183
rect 691 174 695 185
rect 768 187 770 189
rect 772 187 792 189
rect 768 186 792 187
rect 651 157 653 159
rect 651 152 655 157
rect 651 150 653 152
rect 666 173 695 174
rect 666 171 670 173
rect 672 171 695 173
rect 666 170 695 171
rect 666 164 680 166
rect 682 164 687 166
rect 666 162 687 164
rect 683 156 687 162
rect 683 154 684 156
rect 686 154 687 156
rect 683 153 687 154
rect 691 165 695 170
rect 715 182 720 183
rect 715 180 716 182
rect 718 180 720 182
rect 715 174 720 180
rect 691 163 696 165
rect 691 161 693 163
rect 695 161 696 163
rect 691 156 696 161
rect 691 154 693 156
rect 695 154 696 156
rect 706 173 720 174
rect 706 171 710 173
rect 712 171 720 173
rect 706 170 720 171
rect 740 182 753 183
rect 740 180 743 182
rect 745 180 753 182
rect 740 178 753 180
rect 788 182 792 186
rect 740 177 750 178
rect 748 176 750 177
rect 752 176 753 178
rect 732 166 737 167
rect 714 165 727 166
rect 731 165 737 166
rect 714 163 720 165
rect 722 163 734 165
rect 736 163 737 165
rect 714 162 737 163
rect 723 160 737 162
rect 748 169 753 176
rect 788 180 789 182
rect 791 180 792 182
rect 691 152 696 154
rect 651 146 664 150
rect 651 145 655 146
rect 723 153 727 160
rect 732 151 737 160
rect 732 145 744 151
rect 788 158 792 180
rect 776 156 792 158
rect 776 154 778 156
rect 780 154 792 156
rect 776 153 792 154
rect 796 187 808 191
rect 796 185 798 187
rect 800 185 808 187
rect 873 189 897 190
rect 796 165 800 185
rect 873 187 875 189
rect 877 187 897 189
rect 873 186 897 187
rect 820 182 825 183
rect 820 180 821 182
rect 823 180 825 182
rect 820 174 825 180
rect 796 163 801 165
rect 796 161 798 163
rect 800 161 801 163
rect 796 156 801 161
rect 796 154 798 156
rect 800 154 801 156
rect 811 173 825 174
rect 811 171 815 173
rect 817 171 825 173
rect 811 170 825 171
rect 845 182 858 183
rect 845 180 848 182
rect 850 180 858 182
rect 845 178 858 180
rect 845 177 855 178
rect 853 176 855 177
rect 857 176 858 178
rect 837 166 842 167
rect 819 165 832 166
rect 836 165 842 166
rect 819 163 825 165
rect 827 164 839 165
rect 827 163 833 164
rect 819 162 833 163
rect 835 163 839 164
rect 841 163 842 165
rect 835 162 842 163
rect 828 160 842 162
rect 853 169 858 176
rect 796 152 801 154
rect 828 153 832 160
rect 837 151 842 160
rect 837 145 849 151
rect 893 158 897 186
rect 941 187 953 191
rect 941 185 943 187
rect 945 185 953 187
rect 1018 189 1042 190
rect 881 156 897 158
rect 881 154 883 156
rect 885 154 897 156
rect 881 153 897 154
rect 901 182 906 184
rect 901 180 903 182
rect 905 180 906 182
rect 901 178 906 180
rect 901 164 905 178
rect 901 162 902 164
rect 904 162 905 164
rect 901 159 905 162
rect 933 174 937 183
rect 941 174 945 185
rect 1018 187 1020 189
rect 1022 187 1042 189
rect 1018 186 1042 187
rect 901 157 903 159
rect 901 152 905 157
rect 901 150 903 152
rect 916 173 945 174
rect 916 171 920 173
rect 922 171 945 173
rect 916 170 945 171
rect 916 164 930 166
rect 932 164 937 166
rect 916 162 937 164
rect 933 156 937 162
rect 933 154 934 156
rect 936 154 937 156
rect 933 153 937 154
rect 941 165 945 170
rect 965 182 970 183
rect 965 180 966 182
rect 968 180 970 182
rect 965 174 970 180
rect 941 163 946 165
rect 941 161 943 163
rect 945 161 946 163
rect 941 156 946 161
rect 941 154 943 156
rect 945 154 946 156
rect 956 173 970 174
rect 956 171 960 173
rect 962 171 970 173
rect 956 170 970 171
rect 990 182 1003 183
rect 990 180 993 182
rect 995 180 1003 182
rect 990 178 1003 180
rect 1038 182 1042 186
rect 990 177 1000 178
rect 998 176 1000 177
rect 1002 176 1003 178
rect 982 166 987 167
rect 964 165 977 166
rect 981 165 987 166
rect 964 163 970 165
rect 972 163 984 165
rect 986 163 987 165
rect 964 162 987 163
rect 973 160 987 162
rect 998 169 1003 176
rect 1038 180 1039 182
rect 1041 180 1042 182
rect 941 152 946 154
rect 901 146 914 150
rect 901 145 905 146
rect 973 153 977 160
rect 982 151 987 160
rect 982 145 994 151
rect 1038 158 1042 180
rect 1026 156 1042 158
rect 1026 154 1028 156
rect 1030 154 1042 156
rect 1026 153 1042 154
rect 1046 187 1058 191
rect 1046 185 1048 187
rect 1050 185 1058 187
rect 1123 189 1147 190
rect 1046 165 1050 185
rect 1123 187 1125 189
rect 1127 187 1147 189
rect 1123 186 1147 187
rect 1070 182 1075 183
rect 1070 180 1071 182
rect 1073 180 1075 182
rect 1070 174 1075 180
rect 1046 163 1051 165
rect 1046 161 1048 163
rect 1050 161 1051 163
rect 1046 156 1051 161
rect 1046 154 1048 156
rect 1050 154 1051 156
rect 1061 173 1075 174
rect 1061 171 1065 173
rect 1067 171 1075 173
rect 1061 170 1075 171
rect 1095 182 1108 183
rect 1095 180 1098 182
rect 1100 180 1108 182
rect 1095 178 1108 180
rect 1095 177 1105 178
rect 1103 176 1105 177
rect 1107 176 1108 178
rect 1087 166 1092 167
rect 1069 165 1082 166
rect 1086 165 1092 166
rect 1069 163 1075 165
rect 1077 163 1089 165
rect 1091 163 1092 165
rect 1069 162 1092 163
rect 1078 160 1092 162
rect 1103 169 1108 176
rect 1046 152 1051 154
rect 1078 153 1082 160
rect 1087 151 1092 160
rect 1087 145 1099 151
rect 1143 158 1147 186
rect 1131 156 1147 158
rect 1131 154 1133 156
rect 1135 154 1147 156
rect 1131 153 1147 154
rect 147 139 1151 140
rect 147 137 154 139
rect 156 137 194 139
rect 196 137 268 139
rect 270 137 299 139
rect 301 137 373 139
rect 375 137 404 139
rect 406 137 444 139
rect 446 137 518 139
rect 520 137 549 139
rect 551 137 623 139
rect 625 137 654 139
rect 656 137 694 139
rect 696 137 768 139
rect 770 137 799 139
rect 801 137 873 139
rect 875 137 904 139
rect 906 137 944 139
rect 946 137 1018 139
rect 1020 137 1049 139
rect 1051 137 1123 139
rect 1125 137 1151 139
rect 147 132 1151 137
rect 146 127 1150 132
rect 146 125 153 127
rect 155 125 193 127
rect 195 125 267 127
rect 269 125 298 127
rect 300 125 372 127
rect 374 125 403 127
rect 405 125 443 127
rect 445 125 517 127
rect 519 125 548 127
rect 550 125 622 127
rect 624 125 653 127
rect 655 125 693 127
rect 695 125 767 127
rect 769 125 798 127
rect 800 125 872 127
rect 874 125 903 127
rect 905 125 943 127
rect 945 125 1017 127
rect 1019 125 1048 127
rect 1050 125 1122 127
rect 1124 125 1150 127
rect 146 124 1150 125
rect 150 118 154 119
rect 150 114 163 118
rect 150 112 152 114
rect 150 107 154 112
rect 150 105 152 107
rect 150 86 154 105
rect 182 110 186 111
rect 182 108 183 110
rect 185 108 186 110
rect 182 102 186 108
rect 165 100 186 102
rect 165 98 179 100
rect 181 98 186 100
rect 190 110 195 112
rect 190 108 192 110
rect 194 108 195 110
rect 231 113 243 119
rect 190 103 195 108
rect 190 101 192 103
rect 194 101 195 103
rect 190 99 195 101
rect 190 94 194 99
rect 150 84 155 86
rect 150 82 152 84
rect 154 82 155 84
rect 150 80 155 82
rect 165 93 194 94
rect 165 91 169 93
rect 171 91 194 93
rect 165 90 194 91
rect 182 81 186 90
rect 190 79 194 90
rect 222 104 226 111
rect 231 104 236 113
rect 222 102 236 104
rect 213 101 236 102
rect 213 99 219 101
rect 221 99 233 101
rect 235 99 236 101
rect 213 98 226 99
rect 230 98 236 99
rect 231 97 236 98
rect 205 93 219 94
rect 205 91 209 93
rect 211 91 219 93
rect 205 90 219 91
rect 190 77 192 79
rect 194 77 202 79
rect 190 73 202 77
rect 214 84 219 90
rect 214 82 215 84
rect 217 82 219 84
rect 214 81 219 82
rect 247 88 252 95
rect 275 110 291 111
rect 275 108 277 110
rect 279 108 291 110
rect 275 106 291 108
rect 247 87 249 88
rect 239 86 249 87
rect 251 86 252 88
rect 239 84 252 86
rect 239 82 242 84
rect 244 82 252 84
rect 239 81 252 82
rect 287 84 291 106
rect 287 82 288 84
rect 290 82 291 84
rect 287 78 291 82
rect 267 77 291 78
rect 267 75 269 77
rect 271 75 291 77
rect 267 74 291 75
rect 295 110 300 112
rect 295 108 297 110
rect 299 108 300 110
rect 336 113 348 119
rect 400 118 404 119
rect 295 103 300 108
rect 295 101 297 103
rect 299 101 300 103
rect 295 99 300 101
rect 295 79 299 99
rect 327 104 331 111
rect 336 104 341 113
rect 400 114 413 118
rect 400 112 402 114
rect 327 102 341 104
rect 318 101 330 102
rect 318 99 324 101
rect 326 100 330 101
rect 332 101 341 102
rect 332 100 338 101
rect 326 99 338 100
rect 340 99 341 101
rect 318 98 331 99
rect 335 98 341 99
rect 336 97 341 98
rect 310 93 324 94
rect 310 91 314 93
rect 316 91 324 93
rect 310 90 324 91
rect 295 77 297 79
rect 299 77 307 79
rect 295 73 307 77
rect 319 84 324 90
rect 319 82 320 84
rect 322 82 324 84
rect 319 81 324 82
rect 352 88 357 95
rect 380 110 396 111
rect 380 108 382 110
rect 384 108 396 110
rect 380 106 396 108
rect 352 87 354 88
rect 344 86 354 87
rect 356 86 357 88
rect 344 84 357 86
rect 344 82 347 84
rect 349 82 357 84
rect 344 81 357 82
rect 392 78 396 106
rect 400 107 404 112
rect 400 105 402 107
rect 400 102 404 105
rect 432 110 436 111
rect 432 108 433 110
rect 435 108 436 110
rect 400 100 401 102
rect 403 100 404 102
rect 400 86 404 100
rect 432 102 436 108
rect 415 100 436 102
rect 415 98 429 100
rect 431 98 436 100
rect 440 110 445 112
rect 440 108 442 110
rect 444 108 445 110
rect 481 113 493 119
rect 440 103 445 108
rect 440 101 442 103
rect 444 101 445 103
rect 440 99 445 101
rect 440 94 444 99
rect 400 84 405 86
rect 400 82 402 84
rect 404 82 405 84
rect 400 80 405 82
rect 415 93 444 94
rect 415 91 419 93
rect 421 91 444 93
rect 415 90 444 91
rect 432 81 436 90
rect 372 77 396 78
rect 372 75 374 77
rect 376 75 396 77
rect 372 74 396 75
rect 440 79 444 90
rect 472 104 476 111
rect 481 104 486 113
rect 472 102 486 104
rect 463 101 486 102
rect 463 99 469 101
rect 471 99 483 101
rect 485 99 486 101
rect 463 98 476 99
rect 480 98 486 99
rect 481 97 486 98
rect 455 93 469 94
rect 455 91 459 93
rect 461 91 469 93
rect 455 90 469 91
rect 440 77 442 79
rect 444 77 452 79
rect 440 73 452 77
rect 464 84 469 90
rect 464 82 465 84
rect 467 82 469 84
rect 464 81 469 82
rect 497 88 502 95
rect 525 110 541 111
rect 525 108 527 110
rect 529 108 541 110
rect 525 106 541 108
rect 497 87 499 88
rect 489 86 499 87
rect 501 86 502 88
rect 489 84 502 86
rect 489 82 492 84
rect 494 82 502 84
rect 489 81 502 82
rect 537 84 541 106
rect 537 82 538 84
rect 540 82 541 84
rect 537 78 541 82
rect 517 77 541 78
rect 517 75 519 77
rect 521 75 541 77
rect 517 74 541 75
rect 545 110 550 112
rect 545 108 547 110
rect 549 108 550 110
rect 586 113 598 119
rect 650 118 654 119
rect 545 103 550 108
rect 545 101 547 103
rect 549 101 550 103
rect 545 99 550 101
rect 545 79 549 99
rect 577 104 581 111
rect 586 104 591 113
rect 650 114 663 118
rect 650 112 652 114
rect 577 102 591 104
rect 568 101 582 102
rect 568 99 574 101
rect 576 100 582 101
rect 584 101 591 102
rect 584 100 588 101
rect 576 99 588 100
rect 590 99 591 101
rect 568 98 581 99
rect 585 98 591 99
rect 586 97 591 98
rect 560 93 574 94
rect 560 91 564 93
rect 566 91 574 93
rect 560 90 574 91
rect 545 77 547 79
rect 549 77 557 79
rect 545 73 557 77
rect 569 84 574 90
rect 569 82 570 84
rect 572 82 574 84
rect 569 81 574 82
rect 602 88 607 95
rect 630 110 646 111
rect 630 108 632 110
rect 634 108 646 110
rect 630 106 646 108
rect 602 87 604 88
rect 594 86 604 87
rect 606 86 607 88
rect 594 84 607 86
rect 594 82 597 84
rect 599 82 607 84
rect 594 81 607 82
rect 642 78 646 106
rect 650 107 654 112
rect 650 105 652 107
rect 650 102 654 105
rect 682 110 686 111
rect 682 108 683 110
rect 685 108 686 110
rect 650 100 651 102
rect 653 100 654 102
rect 650 86 654 100
rect 682 102 686 108
rect 665 100 686 102
rect 665 98 679 100
rect 681 98 686 100
rect 690 110 695 112
rect 690 108 692 110
rect 694 108 695 110
rect 731 113 743 119
rect 690 103 695 108
rect 690 101 692 103
rect 694 101 695 103
rect 690 99 695 101
rect 690 94 694 99
rect 650 84 655 86
rect 650 82 652 84
rect 654 82 655 84
rect 650 80 655 82
rect 665 93 694 94
rect 665 91 669 93
rect 671 91 694 93
rect 665 90 694 91
rect 682 81 686 90
rect 622 77 646 78
rect 622 75 624 77
rect 626 75 646 77
rect 622 74 646 75
rect 690 79 694 90
rect 722 104 726 111
rect 731 104 736 113
rect 722 102 736 104
rect 713 101 736 102
rect 713 99 719 101
rect 721 99 733 101
rect 735 99 736 101
rect 713 98 726 99
rect 730 98 736 99
rect 731 97 736 98
rect 705 93 719 94
rect 705 91 709 93
rect 711 91 719 93
rect 705 90 719 91
rect 690 77 692 79
rect 694 77 702 79
rect 690 73 702 77
rect 714 84 719 90
rect 714 82 715 84
rect 717 82 719 84
rect 714 81 719 82
rect 747 88 752 95
rect 775 110 791 111
rect 775 108 777 110
rect 779 108 791 110
rect 775 106 791 108
rect 747 87 749 88
rect 739 86 749 87
rect 751 86 752 88
rect 739 84 752 86
rect 739 82 742 84
rect 744 82 752 84
rect 739 81 752 82
rect 787 84 791 106
rect 787 82 788 84
rect 790 82 791 84
rect 787 78 791 82
rect 767 77 791 78
rect 767 75 769 77
rect 771 75 791 77
rect 767 74 791 75
rect 795 110 800 112
rect 795 108 797 110
rect 799 108 800 110
rect 836 113 848 119
rect 900 118 904 119
rect 795 103 800 108
rect 795 101 797 103
rect 799 101 800 103
rect 795 99 800 101
rect 795 79 799 99
rect 827 104 831 111
rect 836 104 841 113
rect 900 114 913 118
rect 900 112 902 114
rect 827 102 841 104
rect 818 101 832 102
rect 818 99 824 101
rect 826 100 832 101
rect 834 101 841 102
rect 834 100 838 101
rect 826 99 838 100
rect 840 99 841 101
rect 818 98 831 99
rect 835 98 841 99
rect 836 97 841 98
rect 810 93 824 94
rect 810 91 814 93
rect 816 91 824 93
rect 810 90 824 91
rect 795 77 797 79
rect 799 77 807 79
rect 795 73 807 77
rect 819 84 824 90
rect 819 82 820 84
rect 822 82 824 84
rect 819 81 824 82
rect 852 88 857 95
rect 880 110 896 111
rect 880 108 882 110
rect 884 108 896 110
rect 880 106 896 108
rect 852 87 854 88
rect 844 86 854 87
rect 856 86 857 88
rect 844 84 857 86
rect 844 82 847 84
rect 849 82 857 84
rect 844 81 857 82
rect 892 78 896 106
rect 900 107 904 112
rect 900 105 902 107
rect 900 102 904 105
rect 932 110 936 111
rect 932 108 933 110
rect 935 108 936 110
rect 900 100 901 102
rect 903 100 904 102
rect 900 86 904 100
rect 932 102 936 108
rect 915 100 936 102
rect 915 98 929 100
rect 931 98 936 100
rect 940 110 945 112
rect 940 108 942 110
rect 944 108 945 110
rect 981 113 993 119
rect 940 103 945 108
rect 940 101 942 103
rect 944 101 945 103
rect 940 99 945 101
rect 940 94 944 99
rect 900 84 905 86
rect 900 82 902 84
rect 904 82 905 84
rect 900 80 905 82
rect 915 93 944 94
rect 915 91 919 93
rect 921 91 944 93
rect 915 90 944 91
rect 932 81 936 90
rect 872 77 896 78
rect 872 75 874 77
rect 876 75 896 77
rect 872 74 896 75
rect 940 79 944 90
rect 972 104 976 111
rect 981 104 986 113
rect 972 102 986 104
rect 963 101 986 102
rect 963 99 969 101
rect 971 99 983 101
rect 985 99 986 101
rect 963 98 976 99
rect 980 98 986 99
rect 981 97 986 98
rect 955 93 969 94
rect 955 91 959 93
rect 961 91 969 93
rect 955 90 969 91
rect 940 77 942 79
rect 944 77 952 79
rect 940 73 952 77
rect 964 84 969 90
rect 964 82 965 84
rect 967 82 969 84
rect 964 81 969 82
rect 997 88 1002 95
rect 1025 110 1041 111
rect 1025 108 1027 110
rect 1029 108 1041 110
rect 1025 106 1041 108
rect 997 87 999 88
rect 989 86 999 87
rect 1001 86 1002 88
rect 989 84 1002 86
rect 989 82 992 84
rect 994 82 1002 84
rect 989 81 1002 82
rect 1037 84 1041 106
rect 1037 82 1038 84
rect 1040 82 1041 84
rect 1037 78 1041 82
rect 1017 77 1041 78
rect 1017 75 1019 77
rect 1021 75 1041 77
rect 1017 74 1041 75
rect 1045 110 1050 112
rect 1045 108 1047 110
rect 1049 108 1050 110
rect 1086 113 1098 119
rect 1045 103 1050 108
rect 1045 101 1047 103
rect 1049 101 1050 103
rect 1045 99 1050 101
rect 1045 79 1049 99
rect 1077 104 1081 111
rect 1086 104 1091 113
rect 1077 102 1091 104
rect 1068 101 1091 102
rect 1068 99 1074 101
rect 1076 99 1082 101
rect 1084 99 1088 101
rect 1090 99 1091 101
rect 1068 98 1091 99
rect 1086 97 1091 98
rect 1060 93 1074 94
rect 1060 91 1064 93
rect 1066 91 1074 93
rect 1060 90 1074 91
rect 1045 77 1047 79
rect 1049 77 1057 79
rect 1045 73 1057 77
rect 1069 84 1074 90
rect 1069 82 1070 84
rect 1072 82 1074 84
rect 1069 81 1074 82
rect 1102 88 1107 95
rect 1130 110 1146 111
rect 1130 108 1132 110
rect 1134 108 1146 110
rect 1130 106 1146 108
rect 1102 87 1104 88
rect 1094 86 1104 87
rect 1106 86 1107 88
rect 1094 84 1107 86
rect 1094 82 1097 84
rect 1099 82 1107 84
rect 1094 81 1107 82
rect 1142 78 1146 106
rect 1122 77 1146 78
rect 1122 75 1124 77
rect 1126 75 1146 77
rect 1122 74 1146 75
rect 146 67 1150 68
rect 146 65 153 67
rect 155 65 193 67
rect 195 65 203 67
rect 205 65 234 67
rect 236 66 287 67
rect 236 65 243 66
rect 146 64 243 65
rect 245 65 287 66
rect 289 65 298 67
rect 300 65 308 67
rect 310 65 339 67
rect 341 65 392 67
rect 394 65 403 67
rect 405 65 443 67
rect 445 65 453 67
rect 455 65 484 67
rect 486 65 493 67
rect 495 65 537 67
rect 539 65 548 67
rect 550 65 558 67
rect 560 65 589 67
rect 591 65 642 67
rect 644 65 653 67
rect 655 65 693 67
rect 695 65 703 67
rect 705 65 734 67
rect 736 65 787 67
rect 789 65 798 67
rect 800 65 808 67
rect 810 65 839 67
rect 841 65 892 67
rect 894 65 903 67
rect 905 65 943 67
rect 945 65 953 67
rect 955 65 984 67
rect 986 65 1037 67
rect 1039 65 1048 67
rect 1050 65 1058 67
rect 1060 66 1089 67
rect 1060 65 1082 66
rect 245 64 1082 65
rect 1084 65 1089 66
rect 1091 65 1142 67
rect 1144 65 1150 67
rect 1084 64 1150 65
rect 146 60 1150 64
rect 145 56 1149 60
rect 145 55 1081 56
rect 145 53 152 55
rect 154 53 192 55
rect 194 53 202 55
rect 204 53 233 55
rect 235 53 286 55
rect 288 53 297 55
rect 299 53 307 55
rect 309 53 338 55
rect 340 53 391 55
rect 393 53 402 55
rect 404 53 442 55
rect 444 53 452 55
rect 454 53 483 55
rect 485 53 492 55
rect 494 53 536 55
rect 538 53 547 55
rect 549 53 557 55
rect 559 53 588 55
rect 590 53 641 55
rect 643 53 652 55
rect 654 53 692 55
rect 694 53 702 55
rect 704 53 733 55
rect 735 53 786 55
rect 788 53 797 55
rect 799 53 807 55
rect 809 53 838 55
rect 840 53 891 55
rect 893 53 902 55
rect 904 53 942 55
rect 944 53 952 55
rect 954 53 983 55
rect 985 53 1036 55
rect 1038 53 1047 55
rect 1049 53 1057 55
rect 1059 54 1081 55
rect 1083 55 1149 56
rect 1083 54 1088 55
rect 1059 53 1088 54
rect 1090 53 1141 55
rect 1143 53 1149 55
rect 145 52 1149 53
rect 189 43 201 47
rect 189 41 191 43
rect 193 41 201 43
rect 266 45 290 46
rect 149 38 154 40
rect 149 36 151 38
rect 153 36 154 38
rect 149 34 154 36
rect 149 15 153 34
rect 181 30 185 39
rect 189 30 193 41
rect 266 43 268 45
rect 270 43 290 45
rect 266 42 290 43
rect 149 13 151 15
rect 149 8 153 13
rect 149 6 151 8
rect 164 29 193 30
rect 164 27 168 29
rect 170 27 193 29
rect 164 26 193 27
rect 164 20 178 22
rect 180 20 185 22
rect 164 18 185 20
rect 181 12 185 18
rect 181 10 182 12
rect 184 10 185 12
rect 181 9 185 10
rect 189 21 193 26
rect 213 38 218 39
rect 213 36 214 38
rect 216 36 218 38
rect 213 30 218 36
rect 189 19 194 21
rect 189 17 191 19
rect 193 17 194 19
rect 189 12 194 17
rect 189 10 191 12
rect 193 10 194 12
rect 204 29 218 30
rect 204 27 208 29
rect 210 27 218 29
rect 204 26 218 27
rect 238 38 251 39
rect 238 36 241 38
rect 243 36 251 38
rect 238 34 251 36
rect 286 38 290 42
rect 238 33 248 34
rect 246 32 248 33
rect 250 32 251 34
rect 230 22 235 23
rect 212 21 225 22
rect 229 21 235 22
rect 212 19 218 21
rect 220 19 232 21
rect 234 19 235 21
rect 212 18 235 19
rect 221 16 235 18
rect 246 25 251 32
rect 286 36 287 38
rect 289 36 290 38
rect 189 8 194 10
rect 149 2 162 6
rect 149 1 153 2
rect 221 9 225 16
rect 230 7 235 16
rect 230 1 242 7
rect 286 14 290 36
rect 274 12 290 14
rect 274 10 276 12
rect 278 10 290 12
rect 274 9 290 10
rect 294 43 306 47
rect 294 41 296 43
rect 298 41 306 43
rect 371 45 395 46
rect 294 21 298 41
rect 371 43 373 45
rect 375 43 395 45
rect 371 42 395 43
rect 318 38 323 39
rect 318 36 319 38
rect 321 36 323 38
rect 318 30 323 36
rect 294 19 299 21
rect 294 17 296 19
rect 298 17 299 19
rect 294 12 299 17
rect 294 10 296 12
rect 298 10 299 12
rect 309 29 323 30
rect 309 27 313 29
rect 315 27 323 29
rect 309 26 323 27
rect 343 38 356 39
rect 343 36 346 38
rect 348 36 356 38
rect 343 34 356 36
rect 343 33 353 34
rect 351 32 353 33
rect 355 32 356 34
rect 335 22 340 23
rect 317 21 330 22
rect 334 21 340 22
rect 317 19 323 21
rect 325 20 337 21
rect 325 19 329 20
rect 317 18 329 19
rect 331 19 337 20
rect 339 19 340 21
rect 331 18 340 19
rect 326 16 340 18
rect 351 25 356 32
rect 294 8 299 10
rect 326 9 330 16
rect 335 7 340 16
rect 335 1 347 7
rect 391 14 395 42
rect 439 43 451 47
rect 439 41 441 43
rect 443 41 451 43
rect 516 45 540 46
rect 379 12 395 14
rect 379 10 381 12
rect 383 10 395 12
rect 379 9 395 10
rect 399 38 404 40
rect 399 36 401 38
rect 403 36 404 38
rect 399 34 404 36
rect 399 20 403 34
rect 399 18 400 20
rect 402 18 403 20
rect 399 15 403 18
rect 431 30 435 39
rect 439 30 443 41
rect 516 43 518 45
rect 520 43 540 45
rect 516 42 540 43
rect 399 13 401 15
rect 399 8 403 13
rect 399 6 401 8
rect 414 29 443 30
rect 414 27 418 29
rect 420 27 443 29
rect 414 26 443 27
rect 414 20 428 22
rect 430 20 435 22
rect 414 18 435 20
rect 431 12 435 18
rect 431 10 432 12
rect 434 10 435 12
rect 431 9 435 10
rect 439 21 443 26
rect 463 38 468 39
rect 463 36 464 38
rect 466 36 468 38
rect 463 30 468 36
rect 439 19 444 21
rect 439 17 441 19
rect 443 17 444 19
rect 439 12 444 17
rect 439 10 441 12
rect 443 10 444 12
rect 454 29 468 30
rect 454 27 458 29
rect 460 27 468 29
rect 454 26 468 27
rect 488 38 501 39
rect 488 36 491 38
rect 493 36 501 38
rect 488 34 501 36
rect 536 38 540 42
rect 488 33 498 34
rect 496 32 498 33
rect 500 32 501 34
rect 480 22 485 23
rect 462 21 475 22
rect 479 21 485 22
rect 462 19 468 21
rect 470 19 482 21
rect 484 19 485 21
rect 462 18 485 19
rect 471 16 485 18
rect 496 25 501 32
rect 536 36 537 38
rect 539 36 540 38
rect 439 8 444 10
rect 399 2 412 6
rect 399 1 403 2
rect 471 9 475 16
rect 480 7 485 16
rect 480 1 492 7
rect 536 14 540 36
rect 524 12 540 14
rect 524 10 526 12
rect 528 10 540 12
rect 524 9 540 10
rect 544 43 556 47
rect 544 41 546 43
rect 548 41 556 43
rect 621 45 645 46
rect 544 21 548 41
rect 621 43 623 45
rect 625 43 645 45
rect 621 42 645 43
rect 568 38 573 39
rect 568 36 569 38
rect 571 36 573 38
rect 568 30 573 36
rect 544 19 549 21
rect 544 17 546 19
rect 548 17 549 19
rect 544 12 549 17
rect 544 10 546 12
rect 548 10 549 12
rect 559 29 573 30
rect 559 27 563 29
rect 565 27 573 29
rect 559 26 573 27
rect 593 38 606 39
rect 593 36 596 38
rect 598 36 606 38
rect 593 34 606 36
rect 593 33 603 34
rect 601 32 603 33
rect 605 32 606 34
rect 585 22 590 23
rect 567 21 580 22
rect 584 21 590 22
rect 567 19 573 21
rect 575 20 587 21
rect 575 19 581 20
rect 567 18 581 19
rect 583 19 587 20
rect 589 19 590 21
rect 583 18 590 19
rect 576 16 590 18
rect 601 25 606 32
rect 544 8 549 10
rect 576 9 580 16
rect 585 7 590 16
rect 585 1 597 7
rect 641 14 645 42
rect 689 43 701 47
rect 689 41 691 43
rect 693 41 701 43
rect 766 45 790 46
rect 629 12 645 14
rect 629 10 631 12
rect 633 10 645 12
rect 629 9 645 10
rect 649 38 654 40
rect 649 36 651 38
rect 653 36 654 38
rect 649 34 654 36
rect 649 20 653 34
rect 649 18 650 20
rect 652 18 653 20
rect 649 15 653 18
rect 681 30 685 39
rect 689 30 693 41
rect 766 43 768 45
rect 770 43 790 45
rect 766 42 790 43
rect 649 13 651 15
rect 649 8 653 13
rect 649 6 651 8
rect 664 29 693 30
rect 664 27 668 29
rect 670 27 693 29
rect 664 26 693 27
rect 664 20 678 22
rect 680 20 685 22
rect 664 18 685 20
rect 681 12 685 18
rect 681 10 682 12
rect 684 10 685 12
rect 681 9 685 10
rect 689 21 693 26
rect 713 38 718 39
rect 713 36 714 38
rect 716 36 718 38
rect 713 30 718 36
rect 689 19 694 21
rect 689 17 691 19
rect 693 17 694 19
rect 689 12 694 17
rect 689 10 691 12
rect 693 10 694 12
rect 704 29 718 30
rect 704 27 708 29
rect 710 27 718 29
rect 704 26 718 27
rect 738 38 751 39
rect 738 36 741 38
rect 743 36 751 38
rect 738 34 751 36
rect 786 38 790 42
rect 738 33 748 34
rect 746 32 748 33
rect 750 32 751 34
rect 730 22 735 23
rect 712 21 725 22
rect 729 21 735 22
rect 712 19 718 21
rect 720 19 732 21
rect 734 19 735 21
rect 712 18 735 19
rect 721 16 735 18
rect 746 25 751 32
rect 786 36 787 38
rect 789 36 790 38
rect 689 8 694 10
rect 649 2 662 6
rect 649 1 653 2
rect 721 9 725 16
rect 730 7 735 16
rect 730 1 742 7
rect 786 14 790 36
rect 774 12 790 14
rect 774 10 776 12
rect 778 10 790 12
rect 774 9 790 10
rect 794 43 806 47
rect 794 41 796 43
rect 798 41 806 43
rect 871 45 895 46
rect 794 21 798 41
rect 871 43 873 45
rect 875 43 895 45
rect 871 42 895 43
rect 818 38 823 39
rect 818 36 819 38
rect 821 36 823 38
rect 818 30 823 36
rect 794 19 799 21
rect 794 17 796 19
rect 798 17 799 19
rect 794 12 799 17
rect 794 10 796 12
rect 798 10 799 12
rect 809 29 823 30
rect 809 27 813 29
rect 815 27 823 29
rect 809 26 823 27
rect 843 38 856 39
rect 843 36 846 38
rect 848 36 856 38
rect 843 34 856 36
rect 843 33 853 34
rect 851 32 853 33
rect 855 32 856 34
rect 835 22 840 23
rect 817 21 830 22
rect 834 21 840 22
rect 817 19 823 21
rect 825 20 837 21
rect 825 19 831 20
rect 817 18 831 19
rect 833 19 837 20
rect 839 19 840 21
rect 833 18 840 19
rect 826 16 840 18
rect 851 25 856 32
rect 794 8 799 10
rect 826 9 830 16
rect 835 7 840 16
rect 835 1 847 7
rect 891 14 895 42
rect 939 43 951 47
rect 939 41 941 43
rect 943 41 951 43
rect 1016 45 1040 46
rect 879 12 895 14
rect 879 10 881 12
rect 883 10 895 12
rect 879 9 895 10
rect 899 38 904 40
rect 899 36 901 38
rect 903 36 904 38
rect 899 34 904 36
rect 899 20 903 34
rect 899 18 900 20
rect 902 18 903 20
rect 899 15 903 18
rect 931 30 935 39
rect 939 30 943 41
rect 1016 43 1018 45
rect 1020 43 1040 45
rect 1016 42 1040 43
rect 899 13 901 15
rect 899 8 903 13
rect 899 6 901 8
rect 914 29 943 30
rect 914 27 918 29
rect 920 27 943 29
rect 914 26 943 27
rect 914 20 928 22
rect 930 20 935 22
rect 914 18 935 20
rect 931 12 935 18
rect 931 10 932 12
rect 934 10 935 12
rect 931 9 935 10
rect 939 21 943 26
rect 963 38 968 39
rect 963 36 964 38
rect 966 36 968 38
rect 963 30 968 36
rect 939 19 944 21
rect 939 17 941 19
rect 943 17 944 19
rect 939 12 944 17
rect 939 10 941 12
rect 943 10 944 12
rect 954 29 968 30
rect 954 27 958 29
rect 960 27 968 29
rect 954 26 968 27
rect 988 38 1001 39
rect 988 36 991 38
rect 993 36 1001 38
rect 988 34 1001 36
rect 1036 38 1040 42
rect 988 33 998 34
rect 996 32 998 33
rect 1000 32 1001 34
rect 980 22 985 23
rect 962 21 975 22
rect 979 21 985 22
rect 962 19 968 21
rect 970 19 982 21
rect 984 19 985 21
rect 962 18 985 19
rect 971 16 985 18
rect 996 25 1001 32
rect 1036 36 1037 38
rect 1039 36 1040 38
rect 939 8 944 10
rect 899 2 912 6
rect 899 1 903 2
rect 971 9 975 16
rect 980 7 985 16
rect 980 1 992 7
rect 1036 14 1040 36
rect 1024 12 1040 14
rect 1024 10 1026 12
rect 1028 10 1040 12
rect 1024 9 1040 10
rect 1044 43 1056 47
rect 1044 41 1046 43
rect 1048 41 1056 43
rect 1121 45 1145 46
rect 1044 21 1048 41
rect 1121 43 1123 45
rect 1125 43 1145 45
rect 1121 42 1145 43
rect 1068 38 1073 39
rect 1068 36 1069 38
rect 1071 36 1073 38
rect 1068 30 1073 36
rect 1044 19 1049 21
rect 1044 17 1046 19
rect 1048 17 1049 19
rect 1044 12 1049 17
rect 1044 10 1046 12
rect 1048 10 1049 12
rect 1059 29 1073 30
rect 1059 27 1063 29
rect 1065 27 1073 29
rect 1059 26 1073 27
rect 1093 38 1106 39
rect 1093 36 1096 38
rect 1098 36 1106 38
rect 1093 34 1106 36
rect 1093 33 1103 34
rect 1101 32 1103 33
rect 1105 32 1106 34
rect 1085 22 1090 23
rect 1067 21 1090 22
rect 1067 19 1073 21
rect 1075 19 1081 21
rect 1083 19 1087 21
rect 1089 19 1090 21
rect 1067 18 1090 19
rect 1076 16 1090 18
rect 1101 25 1106 32
rect 1044 8 1049 10
rect 1076 9 1080 16
rect 1085 7 1090 16
rect 1085 1 1097 7
rect 1141 14 1145 42
rect 1129 12 1145 14
rect 1129 10 1131 12
rect 1133 10 1145 12
rect 1129 9 1145 10
rect 145 -5 1149 -4
rect 145 -7 152 -5
rect 154 -7 192 -5
rect 194 -7 266 -5
rect 268 -7 297 -5
rect 299 -7 371 -5
rect 373 -7 402 -5
rect 404 -7 442 -5
rect 444 -7 516 -5
rect 518 -7 547 -5
rect 549 -7 621 -5
rect 623 -7 652 -5
rect 654 -7 692 -5
rect 694 -7 766 -5
rect 768 -7 797 -5
rect 799 -7 871 -5
rect 873 -7 902 -5
rect 904 -7 942 -5
rect 944 -7 1016 -5
rect 1018 -7 1047 -5
rect 1049 -7 1121 -5
rect 1123 -7 1149 -5
rect 145 -12 1149 -7
<< alu2 >>
rect 233 326 365 327
rect 233 324 234 326
rect 236 324 335 326
rect 337 324 362 326
rect 364 324 365 326
rect 233 323 365 324
rect 449 326 581 327
rect 449 324 450 326
rect 452 324 551 326
rect 553 324 578 326
rect 580 324 581 326
rect 449 323 581 324
rect 654 326 786 327
rect 654 324 655 326
rect 657 324 756 326
rect 758 324 783 326
rect 785 324 786 326
rect 654 323 786 324
rect 873 326 1005 327
rect 873 324 874 326
rect 876 324 975 326
rect 977 324 1002 326
rect 1004 324 1005 326
rect 873 323 1005 324
rect 216 317 222 318
rect 216 315 219 317
rect 221 315 222 317
rect 193 301 205 302
rect 193 299 202 301
rect 204 299 205 301
rect 193 297 205 299
rect 193 224 198 297
rect 216 237 222 315
rect 258 317 262 318
rect 258 315 259 317
rect 261 315 262 317
rect 241 302 245 303
rect 241 300 242 302
rect 244 300 245 302
rect 241 276 245 300
rect 233 272 245 276
rect 233 254 237 272
rect 233 252 234 254
rect 236 252 237 254
rect 233 251 237 252
rect 216 235 217 237
rect 219 235 222 237
rect 216 234 222 235
rect 241 245 245 246
rect 241 243 242 245
rect 244 243 245 245
rect 241 224 245 243
rect 258 237 262 315
rect 385 314 389 318
rect 385 312 386 314
rect 388 312 389 314
rect 272 303 357 304
rect 272 301 273 303
rect 275 301 354 303
rect 356 301 357 303
rect 272 300 357 301
rect 385 277 389 312
rect 432 317 438 318
rect 432 315 435 317
rect 437 315 438 317
rect 329 272 389 277
rect 409 301 421 302
rect 409 299 418 301
rect 420 299 421 301
rect 409 297 421 299
rect 329 261 334 272
rect 329 259 330 261
rect 332 259 334 261
rect 329 257 334 259
rect 258 235 259 237
rect 261 235 262 237
rect 258 234 262 235
rect 273 228 338 229
rect 273 226 274 228
rect 276 226 306 228
rect 308 226 333 228
rect 335 226 338 228
rect 273 225 338 226
rect 273 224 311 225
rect 409 224 414 297
rect 432 237 438 315
rect 474 317 478 318
rect 474 315 475 317
rect 477 315 478 317
rect 457 302 461 303
rect 457 300 458 302
rect 460 300 461 302
rect 457 276 461 300
rect 449 272 461 276
rect 449 254 453 272
rect 449 252 450 254
rect 452 252 453 254
rect 449 251 453 252
rect 432 235 433 237
rect 435 235 438 237
rect 432 234 438 235
rect 457 245 461 246
rect 457 243 458 245
rect 460 243 461 245
rect 457 224 461 243
rect 474 237 478 315
rect 601 314 605 318
rect 601 312 602 314
rect 604 312 605 314
rect 488 303 573 304
rect 488 301 489 303
rect 491 301 570 303
rect 572 301 573 303
rect 488 300 573 301
rect 601 277 605 312
rect 637 317 643 318
rect 637 315 640 317
rect 642 315 643 317
rect 545 272 605 277
rect 614 301 626 302
rect 614 299 623 301
rect 625 299 626 301
rect 614 297 626 299
rect 545 261 550 272
rect 545 259 546 261
rect 548 259 550 261
rect 545 257 550 259
rect 474 235 475 237
rect 477 235 478 237
rect 474 234 478 235
rect 489 228 554 229
rect 489 226 490 228
rect 492 226 522 228
rect 524 226 549 228
rect 551 226 554 228
rect 489 225 554 226
rect 489 224 527 225
rect 614 224 619 297
rect 637 237 643 315
rect 679 317 683 318
rect 679 315 680 317
rect 682 315 683 317
rect 662 302 666 303
rect 662 300 663 302
rect 665 300 666 302
rect 662 276 666 300
rect 654 272 666 276
rect 654 254 658 272
rect 654 252 655 254
rect 657 252 658 254
rect 654 251 658 252
rect 637 235 638 237
rect 640 235 643 237
rect 637 234 643 235
rect 662 245 666 246
rect 662 243 663 245
rect 665 243 666 245
rect 662 224 666 243
rect 679 237 683 315
rect 806 314 810 318
rect 806 312 807 314
rect 809 312 810 314
rect 693 303 778 304
rect 693 301 694 303
rect 696 301 775 303
rect 777 301 778 303
rect 693 300 778 301
rect 806 277 810 312
rect 856 317 862 318
rect 856 315 859 317
rect 861 315 862 317
rect 750 272 810 277
rect 833 301 845 302
rect 833 299 842 301
rect 844 299 845 301
rect 833 297 845 299
rect 750 261 755 272
rect 750 259 751 261
rect 753 259 755 261
rect 750 257 755 259
rect 679 235 680 237
rect 682 235 683 237
rect 679 234 683 235
rect 694 228 759 229
rect 694 226 695 228
rect 697 226 727 228
rect 729 226 754 228
rect 756 226 759 228
rect 694 225 759 226
rect 694 224 732 225
rect 833 224 838 297
rect 856 237 862 315
rect 898 317 902 318
rect 898 315 899 317
rect 901 315 902 317
rect 881 302 885 303
rect 881 300 882 302
rect 884 300 885 302
rect 881 276 885 300
rect 873 272 885 276
rect 873 254 877 272
rect 873 252 874 254
rect 876 252 877 254
rect 873 251 877 252
rect 856 235 857 237
rect 859 235 862 237
rect 856 234 862 235
rect 881 245 885 246
rect 881 243 882 245
rect 884 243 885 245
rect 881 224 885 243
rect 898 237 902 315
rect 1025 314 1029 318
rect 1025 312 1026 314
rect 1028 312 1029 314
rect 912 303 997 304
rect 912 301 913 303
rect 915 301 994 303
rect 996 301 997 303
rect 912 300 997 301
rect 1025 277 1029 312
rect 969 272 1029 277
rect 969 261 974 272
rect 969 259 970 261
rect 972 259 974 261
rect 969 257 974 259
rect 898 235 899 237
rect 901 235 902 237
rect 898 234 902 235
rect 913 228 978 229
rect 913 226 914 228
rect 916 226 946 228
rect 948 226 973 228
rect 975 226 978 228
rect 913 225 978 226
rect 1069 228 1102 229
rect 1069 226 1070 228
rect 1072 226 1097 228
rect 1099 226 1102 228
rect 1069 225 1102 226
rect 913 224 951 225
rect 193 220 245 224
rect 409 220 461 224
rect 614 220 666 224
rect 833 220 885 224
rect 215 182 248 183
rect 215 180 216 182
rect 218 180 243 182
rect 245 180 248 182
rect 215 179 248 180
rect 288 182 353 183
rect 288 180 289 182
rect 291 180 321 182
rect 323 180 348 182
rect 350 180 353 182
rect 288 179 353 180
rect 465 182 498 183
rect 465 180 466 182
rect 468 180 493 182
rect 495 180 498 182
rect 465 179 498 180
rect 538 182 603 183
rect 538 180 539 182
rect 541 180 571 182
rect 573 180 598 182
rect 600 180 603 182
rect 538 179 603 180
rect 715 182 748 183
rect 715 180 716 182
rect 718 180 743 182
rect 745 180 748 182
rect 715 179 748 180
rect 788 182 853 183
rect 788 180 789 182
rect 791 180 821 182
rect 823 180 848 182
rect 850 180 853 182
rect 788 179 853 180
rect 965 182 998 183
rect 965 180 966 182
rect 968 180 993 182
rect 995 180 998 182
rect 965 179 998 180
rect 1038 182 1103 183
rect 1038 180 1039 182
rect 1041 180 1071 182
rect 1073 180 1098 182
rect 1100 180 1103 182
rect 1038 179 1103 180
rect 330 164 405 165
rect 330 162 331 164
rect 333 162 402 164
rect 404 162 405 164
rect 330 161 405 162
rect 582 164 655 165
rect 582 162 583 164
rect 585 162 652 164
rect 654 162 655 164
rect 582 161 655 162
rect 832 164 905 165
rect 832 162 833 164
rect 835 162 902 164
rect 904 162 905 164
rect 832 161 905 162
rect 183 156 301 157
rect 183 154 184 156
rect 186 154 298 156
rect 300 154 301 156
rect 183 153 301 154
rect 433 156 551 157
rect 433 154 434 156
rect 436 154 548 156
rect 550 154 551 156
rect 433 153 551 154
rect 683 156 801 157
rect 683 154 684 156
rect 686 154 798 156
rect 800 154 801 156
rect 683 153 801 154
rect 933 156 1051 157
rect 933 154 934 156
rect 936 154 1048 156
rect 1050 154 1051 156
rect 933 153 1051 154
rect 182 110 300 111
rect 182 108 183 110
rect 185 108 297 110
rect 299 108 300 110
rect 182 107 300 108
rect 432 110 550 111
rect 432 108 433 110
rect 435 108 547 110
rect 549 108 550 110
rect 432 107 550 108
rect 682 110 800 111
rect 682 108 683 110
rect 685 108 797 110
rect 799 108 800 110
rect 682 107 800 108
rect 932 110 1050 111
rect 932 108 933 110
rect 935 108 1047 110
rect 1049 108 1050 110
rect 932 107 1050 108
rect 329 102 404 103
rect 329 100 330 102
rect 332 100 401 102
rect 403 100 404 102
rect 329 99 404 100
rect 581 102 654 103
rect 581 100 582 102
rect 584 100 651 102
rect 653 100 654 102
rect 581 99 654 100
rect 831 102 904 103
rect 831 100 832 102
rect 834 100 901 102
rect 903 100 904 102
rect 831 99 904 100
rect 1081 101 1085 102
rect 1081 99 1082 101
rect 1084 99 1085 101
rect 1081 92 1085 99
rect 1081 90 1082 92
rect 1084 90 1085 92
rect 1081 89 1085 90
rect 214 84 247 85
rect 214 82 215 84
rect 217 82 242 84
rect 244 82 247 84
rect 214 81 247 82
rect 287 84 352 85
rect 287 82 288 84
rect 290 82 320 84
rect 322 82 347 84
rect 349 82 352 84
rect 287 81 352 82
rect 464 84 497 85
rect 464 82 465 84
rect 467 82 492 84
rect 494 82 497 84
rect 464 81 497 82
rect 537 84 602 85
rect 537 82 538 84
rect 540 82 570 84
rect 572 82 597 84
rect 599 82 602 84
rect 537 81 602 82
rect 714 84 747 85
rect 714 82 715 84
rect 717 82 742 84
rect 744 82 747 84
rect 714 81 747 82
rect 787 84 852 85
rect 787 82 788 84
rect 790 82 820 84
rect 822 82 847 84
rect 849 82 852 84
rect 787 81 852 82
rect 964 84 997 85
rect 964 82 965 84
rect 967 82 992 84
rect 994 82 997 84
rect 964 81 997 82
rect 1037 84 1102 85
rect 1037 82 1038 84
rect 1040 82 1070 84
rect 1072 82 1097 84
rect 1099 82 1102 84
rect 1037 81 1102 82
rect 241 66 246 81
rect 241 64 243 66
rect 245 64 246 66
rect 491 67 496 81
rect 491 65 493 67
rect 495 65 496 67
rect 491 64 496 65
rect 1081 76 1085 77
rect 1081 74 1082 76
rect 1084 74 1085 76
rect 1081 66 1085 74
rect 1081 64 1082 66
rect 1084 64 1085 66
rect 241 61 246 64
rect 1081 62 1085 64
rect 1080 56 1084 58
rect 490 55 495 56
rect 490 53 492 55
rect 494 53 495 55
rect 490 39 495 53
rect 1080 54 1081 56
rect 1083 54 1084 56
rect 1080 46 1084 54
rect 1080 44 1081 46
rect 1083 44 1084 46
rect 1080 43 1084 44
rect 213 38 246 39
rect 213 36 214 38
rect 216 36 241 38
rect 243 36 246 38
rect 213 35 246 36
rect 286 38 351 39
rect 286 36 287 38
rect 289 36 319 38
rect 321 36 346 38
rect 348 36 351 38
rect 286 35 351 36
rect 463 38 496 39
rect 463 36 464 38
rect 466 36 491 38
rect 493 36 496 38
rect 463 35 496 36
rect 536 38 601 39
rect 536 36 537 38
rect 539 36 569 38
rect 571 36 596 38
rect 598 36 601 38
rect 536 35 601 36
rect 713 38 746 39
rect 713 36 714 38
rect 716 36 741 38
rect 743 36 746 38
rect 713 35 746 36
rect 786 38 851 39
rect 786 36 787 38
rect 789 36 819 38
rect 821 36 846 38
rect 848 36 851 38
rect 786 35 851 36
rect 963 38 996 39
rect 963 36 964 38
rect 966 36 991 38
rect 993 36 996 38
rect 963 35 996 36
rect 1036 38 1101 39
rect 1036 36 1037 38
rect 1039 36 1069 38
rect 1071 36 1096 38
rect 1098 36 1101 38
rect 1036 35 1101 36
rect 1080 30 1084 31
rect 1080 28 1081 30
rect 1083 28 1084 30
rect 1080 21 1084 28
rect 328 20 403 21
rect 328 18 329 20
rect 331 18 400 20
rect 402 18 403 20
rect 328 17 403 18
rect 580 20 653 21
rect 580 18 581 20
rect 583 18 650 20
rect 652 18 653 20
rect 580 17 653 18
rect 830 20 903 21
rect 830 18 831 20
rect 833 18 900 20
rect 902 18 903 20
rect 1080 19 1081 21
rect 1083 19 1084 21
rect 1080 18 1084 19
rect 830 17 903 18
rect 181 12 299 13
rect 181 10 182 12
rect 184 10 296 12
rect 298 10 299 12
rect 181 9 299 10
rect 431 12 549 13
rect 431 10 432 12
rect 434 10 546 12
rect 548 10 549 12
rect 431 9 549 10
rect 681 12 799 13
rect 681 10 682 12
rect 684 10 796 12
rect 798 10 799 12
rect 681 9 799 10
rect 931 12 1049 13
rect 931 10 932 12
rect 934 10 1046 12
rect 1048 10 1049 12
rect 931 9 1049 10
<< alu3 >>
rect 1081 92 1085 93
rect 1081 90 1082 92
rect 1084 90 1085 92
rect 1081 76 1085 90
rect 1081 74 1082 76
rect 1084 74 1085 76
rect 1081 73 1085 74
rect 1080 46 1084 47
rect 1080 44 1081 46
rect 1083 44 1084 46
rect 1080 30 1084 44
rect 1080 28 1081 30
rect 1083 28 1084 30
rect 1080 27 1084 28
<< ptie >>
rect 230 343 236 345
rect 230 341 232 343
rect 234 341 236 343
rect 230 339 236 341
rect 270 343 276 345
rect 270 341 272 343
rect 274 341 276 343
rect 270 339 276 341
rect 341 343 347 345
rect 341 341 343 343
rect 345 341 347 343
rect 341 339 347 341
rect 382 343 388 345
rect 382 341 384 343
rect 386 341 388 343
rect 382 339 388 341
rect 446 343 452 345
rect 446 341 448 343
rect 450 341 452 343
rect 446 339 452 341
rect 486 343 492 345
rect 486 341 488 343
rect 490 341 492 343
rect 486 339 492 341
rect 557 343 563 345
rect 557 341 559 343
rect 561 341 563 343
rect 557 339 563 341
rect 598 343 604 345
rect 598 341 600 343
rect 602 341 604 343
rect 598 339 604 341
rect 651 343 657 345
rect 651 341 653 343
rect 655 341 657 343
rect 651 339 657 341
rect 691 343 697 345
rect 691 341 693 343
rect 695 341 697 343
rect 691 339 697 341
rect 762 343 768 345
rect 762 341 764 343
rect 766 341 768 343
rect 762 339 768 341
rect 803 343 809 345
rect 803 341 805 343
rect 807 341 809 343
rect 803 339 809 341
rect 870 343 876 345
rect 870 341 872 343
rect 874 341 876 343
rect 870 339 876 341
rect 910 343 916 345
rect 910 341 912 343
rect 914 341 916 343
rect 910 339 916 341
rect 981 343 987 345
rect 981 341 983 343
rect 985 341 987 343
rect 981 339 987 341
rect 1022 343 1028 345
rect 1022 341 1024 343
rect 1026 341 1028 343
rect 1022 339 1028 341
rect 202 211 208 213
rect 202 209 204 211
rect 206 209 208 211
rect 202 207 208 209
rect 270 211 276 213
rect 270 209 272 211
rect 274 209 276 211
rect 270 207 276 209
rect 282 211 288 213
rect 282 209 284 211
rect 286 209 288 211
rect 282 207 288 209
rect 323 211 329 213
rect 323 209 325 211
rect 327 209 329 211
rect 323 207 329 209
rect 418 211 424 213
rect 418 209 420 211
rect 422 209 424 211
rect 418 207 424 209
rect 486 211 492 213
rect 486 209 488 211
rect 490 209 492 211
rect 486 207 492 209
rect 498 211 504 213
rect 498 209 500 211
rect 502 209 504 211
rect 498 207 504 209
rect 539 211 545 213
rect 539 209 541 211
rect 543 209 545 211
rect 539 207 545 209
rect 623 211 629 213
rect 623 209 625 211
rect 627 209 629 211
rect 623 207 629 209
rect 691 211 697 213
rect 691 209 693 211
rect 695 209 697 211
rect 691 207 697 209
rect 703 211 709 213
rect 703 209 705 211
rect 707 209 709 211
rect 703 207 709 209
rect 744 211 750 213
rect 744 209 746 211
rect 748 209 750 211
rect 744 207 750 209
rect 842 211 848 213
rect 842 209 844 211
rect 846 209 848 211
rect 842 207 848 209
rect 910 211 916 213
rect 910 209 912 211
rect 914 209 916 211
rect 910 207 916 209
rect 922 211 928 213
rect 922 209 924 211
rect 926 209 928 211
rect 922 207 928 209
rect 963 211 969 213
rect 963 209 965 211
rect 967 209 969 211
rect 963 207 969 209
rect 1046 211 1052 213
rect 1046 209 1048 211
rect 1050 209 1052 211
rect 1046 207 1052 209
rect 1087 211 1093 213
rect 1087 209 1089 211
rect 1091 209 1093 211
rect 1087 207 1093 209
rect 152 199 158 201
rect 152 197 154 199
rect 156 197 158 199
rect 192 199 198 201
rect 192 197 194 199
rect 196 197 198 199
rect 152 195 158 197
rect 192 195 198 197
rect 233 199 239 201
rect 233 197 235 199
rect 237 197 239 199
rect 233 195 239 197
rect 297 199 303 201
rect 297 197 299 199
rect 301 197 303 199
rect 297 195 303 197
rect 338 199 344 201
rect 338 197 340 199
rect 342 197 344 199
rect 338 195 344 197
rect 402 199 408 201
rect 402 197 404 199
rect 406 197 408 199
rect 442 199 448 201
rect 442 197 444 199
rect 446 197 448 199
rect 402 195 408 197
rect 442 195 448 197
rect 483 199 489 201
rect 483 197 485 199
rect 487 197 489 199
rect 483 195 489 197
rect 547 199 553 201
rect 547 197 549 199
rect 551 197 553 199
rect 547 195 553 197
rect 588 199 594 201
rect 588 197 590 199
rect 592 197 594 199
rect 588 195 594 197
rect 652 199 658 201
rect 652 197 654 199
rect 656 197 658 199
rect 692 199 698 201
rect 692 197 694 199
rect 696 197 698 199
rect 652 195 658 197
rect 692 195 698 197
rect 733 199 739 201
rect 733 197 735 199
rect 737 197 739 199
rect 733 195 739 197
rect 797 199 803 201
rect 797 197 799 199
rect 801 197 803 199
rect 797 195 803 197
rect 838 199 844 201
rect 838 197 840 199
rect 842 197 844 199
rect 838 195 844 197
rect 902 199 908 201
rect 902 197 904 199
rect 906 197 908 199
rect 942 199 948 201
rect 942 197 944 199
rect 946 197 948 199
rect 902 195 908 197
rect 942 195 948 197
rect 983 199 989 201
rect 983 197 985 199
rect 987 197 989 199
rect 983 195 989 197
rect 1047 199 1053 201
rect 1047 197 1049 199
rect 1051 197 1053 199
rect 1047 195 1053 197
rect 1088 199 1094 201
rect 1088 197 1090 199
rect 1092 197 1094 199
rect 1088 195 1094 197
rect 151 67 157 69
rect 191 67 197 69
rect 151 65 153 67
rect 155 65 157 67
rect 151 63 157 65
rect 191 65 193 67
rect 195 65 197 67
rect 191 63 197 65
rect 232 67 238 69
rect 232 65 234 67
rect 236 65 238 67
rect 232 63 238 65
rect 296 67 302 69
rect 296 65 298 67
rect 300 65 302 67
rect 296 63 302 65
rect 337 67 343 69
rect 337 65 339 67
rect 341 65 343 67
rect 337 63 343 65
rect 401 67 407 69
rect 441 67 447 69
rect 401 65 403 67
rect 405 65 407 67
rect 401 63 407 65
rect 441 65 443 67
rect 445 65 447 67
rect 441 63 447 65
rect 482 67 488 69
rect 482 65 484 67
rect 486 65 488 67
rect 482 63 488 65
rect 546 67 552 69
rect 546 65 548 67
rect 550 65 552 67
rect 546 63 552 65
rect 587 67 593 69
rect 587 65 589 67
rect 591 65 593 67
rect 587 63 593 65
rect 651 67 657 69
rect 691 67 697 69
rect 651 65 653 67
rect 655 65 657 67
rect 651 63 657 65
rect 691 65 693 67
rect 695 65 697 67
rect 691 63 697 65
rect 732 67 738 69
rect 732 65 734 67
rect 736 65 738 67
rect 732 63 738 65
rect 796 67 802 69
rect 796 65 798 67
rect 800 65 802 67
rect 796 63 802 65
rect 837 67 843 69
rect 837 65 839 67
rect 841 65 843 67
rect 837 63 843 65
rect 901 67 907 69
rect 941 67 947 69
rect 901 65 903 67
rect 905 65 907 67
rect 901 63 907 65
rect 941 65 943 67
rect 945 65 947 67
rect 941 63 947 65
rect 982 67 988 69
rect 982 65 984 67
rect 986 65 988 67
rect 982 63 988 65
rect 1046 67 1052 69
rect 1046 65 1048 67
rect 1050 65 1052 67
rect 1046 63 1052 65
rect 1087 67 1093 69
rect 1087 65 1089 67
rect 1091 65 1093 67
rect 1087 63 1093 65
rect 150 55 156 57
rect 150 53 152 55
rect 154 53 156 55
rect 190 55 196 57
rect 190 53 192 55
rect 194 53 196 55
rect 150 51 156 53
rect 190 51 196 53
rect 231 55 237 57
rect 231 53 233 55
rect 235 53 237 55
rect 231 51 237 53
rect 295 55 301 57
rect 295 53 297 55
rect 299 53 301 55
rect 295 51 301 53
rect 336 55 342 57
rect 336 53 338 55
rect 340 53 342 55
rect 336 51 342 53
rect 400 55 406 57
rect 400 53 402 55
rect 404 53 406 55
rect 440 55 446 57
rect 440 53 442 55
rect 444 53 446 55
rect 400 51 406 53
rect 440 51 446 53
rect 481 55 487 57
rect 481 53 483 55
rect 485 53 487 55
rect 481 51 487 53
rect 545 55 551 57
rect 545 53 547 55
rect 549 53 551 55
rect 545 51 551 53
rect 586 55 592 57
rect 586 53 588 55
rect 590 53 592 55
rect 586 51 592 53
rect 650 55 656 57
rect 650 53 652 55
rect 654 53 656 55
rect 690 55 696 57
rect 690 53 692 55
rect 694 53 696 55
rect 650 51 656 53
rect 690 51 696 53
rect 731 55 737 57
rect 731 53 733 55
rect 735 53 737 55
rect 731 51 737 53
rect 795 55 801 57
rect 795 53 797 55
rect 799 53 801 55
rect 795 51 801 53
rect 836 55 842 57
rect 836 53 838 55
rect 840 53 842 55
rect 836 51 842 53
rect 900 55 906 57
rect 900 53 902 55
rect 904 53 906 55
rect 940 55 946 57
rect 940 53 942 55
rect 944 53 946 55
rect 900 51 906 53
rect 940 51 946 53
rect 981 55 987 57
rect 981 53 983 55
rect 985 53 987 55
rect 981 51 987 53
rect 1045 55 1051 57
rect 1045 53 1047 55
rect 1049 53 1051 55
rect 1045 51 1051 53
rect 1086 55 1092 57
rect 1086 53 1088 55
rect 1090 53 1092 55
rect 1086 51 1092 53
<< ntie >>
rect 230 283 236 285
rect 230 281 232 283
rect 234 281 236 283
rect 230 279 236 281
rect 270 283 276 285
rect 270 281 272 283
rect 274 281 276 283
rect 308 283 314 285
rect 270 279 276 281
rect 308 281 310 283
rect 312 281 314 283
rect 382 283 388 285
rect 308 279 314 281
rect 382 281 384 283
rect 386 281 388 283
rect 382 279 388 281
rect 446 283 452 285
rect 446 281 448 283
rect 450 281 452 283
rect 446 279 452 281
rect 486 283 492 285
rect 486 281 488 283
rect 490 281 492 283
rect 524 283 530 285
rect 486 279 492 281
rect 524 281 526 283
rect 528 281 530 283
rect 598 283 604 285
rect 524 279 530 281
rect 598 281 600 283
rect 602 281 604 283
rect 598 279 604 281
rect 651 283 657 285
rect 651 281 653 283
rect 655 281 657 283
rect 651 279 657 281
rect 691 283 697 285
rect 691 281 693 283
rect 695 281 697 283
rect 729 283 735 285
rect 691 279 697 281
rect 729 281 731 283
rect 733 281 735 283
rect 803 283 809 285
rect 729 279 735 281
rect 803 281 805 283
rect 807 281 809 283
rect 803 279 809 281
rect 870 283 876 285
rect 870 281 872 283
rect 874 281 876 283
rect 870 279 876 281
rect 910 283 916 285
rect 910 281 912 283
rect 914 281 916 283
rect 948 283 954 285
rect 910 279 916 281
rect 948 281 950 283
rect 952 281 954 283
rect 1022 283 1028 285
rect 948 279 954 281
rect 1022 281 1024 283
rect 1026 281 1028 283
rect 1022 279 1028 281
rect 202 271 208 273
rect 202 269 204 271
rect 206 269 208 271
rect 202 267 208 269
rect 270 271 276 273
rect 270 269 272 271
rect 274 269 276 271
rect 270 267 276 269
rect 282 271 288 273
rect 282 269 284 271
rect 286 269 288 271
rect 356 271 362 273
rect 282 267 288 269
rect 356 269 358 271
rect 360 269 362 271
rect 418 271 424 273
rect 356 267 362 269
rect 418 269 420 271
rect 422 269 424 271
rect 418 267 424 269
rect 486 271 492 273
rect 486 269 488 271
rect 490 269 492 271
rect 486 267 492 269
rect 498 271 504 273
rect 498 269 500 271
rect 502 269 504 271
rect 572 271 578 273
rect 498 267 504 269
rect 572 269 574 271
rect 576 269 578 271
rect 623 271 629 273
rect 572 267 578 269
rect 623 269 625 271
rect 627 269 629 271
rect 623 267 629 269
rect 691 271 697 273
rect 691 269 693 271
rect 695 269 697 271
rect 691 267 697 269
rect 703 271 709 273
rect 703 269 705 271
rect 707 269 709 271
rect 777 271 783 273
rect 703 267 709 269
rect 777 269 779 271
rect 781 269 783 271
rect 842 271 848 273
rect 777 267 783 269
rect 842 269 844 271
rect 846 269 848 271
rect 842 267 848 269
rect 910 271 916 273
rect 910 269 912 271
rect 914 269 916 271
rect 910 267 916 269
rect 922 271 928 273
rect 922 269 924 271
rect 926 269 928 271
rect 996 271 1002 273
rect 922 267 928 269
rect 996 269 998 271
rect 1000 269 1002 271
rect 1046 271 1052 273
rect 996 267 1002 269
rect 1046 269 1048 271
rect 1050 269 1052 271
rect 1120 271 1126 273
rect 1046 267 1052 269
rect 1120 269 1122 271
rect 1124 269 1126 271
rect 1120 267 1126 269
rect 152 139 158 141
rect 152 137 154 139
rect 156 137 158 139
rect 192 139 198 141
rect 152 135 158 137
rect 192 137 194 139
rect 196 137 198 139
rect 266 139 272 141
rect 192 135 198 137
rect 266 137 268 139
rect 270 137 272 139
rect 297 139 303 141
rect 266 135 272 137
rect 297 137 299 139
rect 301 137 303 139
rect 371 139 377 141
rect 297 135 303 137
rect 371 137 373 139
rect 375 137 377 139
rect 402 139 408 141
rect 371 135 377 137
rect 402 137 404 139
rect 406 137 408 139
rect 442 139 448 141
rect 402 135 408 137
rect 442 137 444 139
rect 446 137 448 139
rect 516 139 522 141
rect 442 135 448 137
rect 516 137 518 139
rect 520 137 522 139
rect 547 139 553 141
rect 516 135 522 137
rect 547 137 549 139
rect 551 137 553 139
rect 621 139 627 141
rect 547 135 553 137
rect 621 137 623 139
rect 625 137 627 139
rect 652 139 658 141
rect 621 135 627 137
rect 652 137 654 139
rect 656 137 658 139
rect 692 139 698 141
rect 652 135 658 137
rect 692 137 694 139
rect 696 137 698 139
rect 766 139 772 141
rect 692 135 698 137
rect 766 137 768 139
rect 770 137 772 139
rect 797 139 803 141
rect 766 135 772 137
rect 797 137 799 139
rect 801 137 803 139
rect 871 139 877 141
rect 797 135 803 137
rect 871 137 873 139
rect 875 137 877 139
rect 902 139 908 141
rect 871 135 877 137
rect 902 137 904 139
rect 906 137 908 139
rect 942 139 948 141
rect 902 135 908 137
rect 942 137 944 139
rect 946 137 948 139
rect 1016 139 1022 141
rect 942 135 948 137
rect 1016 137 1018 139
rect 1020 137 1022 139
rect 1047 139 1053 141
rect 1016 135 1022 137
rect 1047 137 1049 139
rect 1051 137 1053 139
rect 1121 139 1127 141
rect 1047 135 1053 137
rect 1121 137 1123 139
rect 1125 137 1127 139
rect 1121 135 1127 137
rect 151 127 157 129
rect 151 125 153 127
rect 155 125 157 127
rect 191 127 197 129
rect 151 123 157 125
rect 191 125 193 127
rect 195 125 197 127
rect 265 127 271 129
rect 191 123 197 125
rect 265 125 267 127
rect 269 125 271 127
rect 296 127 302 129
rect 265 123 271 125
rect 296 125 298 127
rect 300 125 302 127
rect 370 127 376 129
rect 296 123 302 125
rect 370 125 372 127
rect 374 125 376 127
rect 401 127 407 129
rect 370 123 376 125
rect 401 125 403 127
rect 405 125 407 127
rect 441 127 447 129
rect 401 123 407 125
rect 441 125 443 127
rect 445 125 447 127
rect 515 127 521 129
rect 441 123 447 125
rect 515 125 517 127
rect 519 125 521 127
rect 546 127 552 129
rect 515 123 521 125
rect 546 125 548 127
rect 550 125 552 127
rect 620 127 626 129
rect 546 123 552 125
rect 620 125 622 127
rect 624 125 626 127
rect 651 127 657 129
rect 620 123 626 125
rect 651 125 653 127
rect 655 125 657 127
rect 691 127 697 129
rect 651 123 657 125
rect 691 125 693 127
rect 695 125 697 127
rect 765 127 771 129
rect 691 123 697 125
rect 765 125 767 127
rect 769 125 771 127
rect 796 127 802 129
rect 765 123 771 125
rect 796 125 798 127
rect 800 125 802 127
rect 870 127 876 129
rect 796 123 802 125
rect 870 125 872 127
rect 874 125 876 127
rect 901 127 907 129
rect 870 123 876 125
rect 901 125 903 127
rect 905 125 907 127
rect 941 127 947 129
rect 901 123 907 125
rect 941 125 943 127
rect 945 125 947 127
rect 1015 127 1021 129
rect 941 123 947 125
rect 1015 125 1017 127
rect 1019 125 1021 127
rect 1046 127 1052 129
rect 1015 123 1021 125
rect 1046 125 1048 127
rect 1050 125 1052 127
rect 1120 127 1126 129
rect 1046 123 1052 125
rect 1120 125 1122 127
rect 1124 125 1126 127
rect 1120 123 1126 125
rect 150 -5 156 -3
rect 150 -7 152 -5
rect 154 -7 156 -5
rect 190 -5 196 -3
rect 150 -9 156 -7
rect 190 -7 192 -5
rect 194 -7 196 -5
rect 264 -5 270 -3
rect 190 -9 196 -7
rect 264 -7 266 -5
rect 268 -7 270 -5
rect 295 -5 301 -3
rect 264 -9 270 -7
rect 295 -7 297 -5
rect 299 -7 301 -5
rect 369 -5 375 -3
rect 295 -9 301 -7
rect 369 -7 371 -5
rect 373 -7 375 -5
rect 400 -5 406 -3
rect 369 -9 375 -7
rect 400 -7 402 -5
rect 404 -7 406 -5
rect 440 -5 446 -3
rect 400 -9 406 -7
rect 440 -7 442 -5
rect 444 -7 446 -5
rect 514 -5 520 -3
rect 440 -9 446 -7
rect 514 -7 516 -5
rect 518 -7 520 -5
rect 545 -5 551 -3
rect 514 -9 520 -7
rect 545 -7 547 -5
rect 549 -7 551 -5
rect 619 -5 625 -3
rect 545 -9 551 -7
rect 619 -7 621 -5
rect 623 -7 625 -5
rect 650 -5 656 -3
rect 619 -9 625 -7
rect 650 -7 652 -5
rect 654 -7 656 -5
rect 690 -5 696 -3
rect 650 -9 656 -7
rect 690 -7 692 -5
rect 694 -7 696 -5
rect 764 -5 770 -3
rect 690 -9 696 -7
rect 764 -7 766 -5
rect 768 -7 770 -5
rect 795 -5 801 -3
rect 764 -9 770 -7
rect 795 -7 797 -5
rect 799 -7 801 -5
rect 869 -5 875 -3
rect 795 -9 801 -7
rect 869 -7 871 -5
rect 873 -7 875 -5
rect 900 -5 906 -3
rect 869 -9 875 -7
rect 900 -7 902 -5
rect 904 -7 906 -5
rect 940 -5 946 -3
rect 900 -9 906 -7
rect 940 -7 942 -5
rect 944 -7 946 -5
rect 1014 -5 1020 -3
rect 940 -9 946 -7
rect 1014 -7 1016 -5
rect 1018 -7 1020 -5
rect 1045 -5 1051 -3
rect 1014 -9 1020 -7
rect 1045 -7 1047 -5
rect 1049 -7 1051 -5
rect 1119 -5 1125 -3
rect 1045 -9 1051 -7
rect 1119 -7 1121 -5
rect 1123 -7 1125 -5
rect 1119 -9 1125 -7
<< nmos >>
rect 208 324 210 335
rect 215 324 217 335
rect 228 324 230 333
rect 248 324 250 335
rect 255 324 257 335
rect 268 324 270 333
rect 296 327 298 339
rect 303 327 305 339
rect 313 327 315 336
rect 323 327 325 336
rect 339 322 341 331
rect 360 324 362 335
rect 367 324 369 335
rect 380 324 382 333
rect 424 324 426 335
rect 431 324 433 335
rect 444 324 446 333
rect 464 324 466 335
rect 471 324 473 335
rect 484 324 486 333
rect 512 327 514 339
rect 519 327 521 339
rect 529 327 531 336
rect 539 327 541 336
rect 555 322 557 331
rect 576 324 578 335
rect 583 324 585 335
rect 596 324 598 333
rect 629 324 631 335
rect 636 324 638 335
rect 649 324 651 333
rect 669 324 671 335
rect 676 324 678 335
rect 689 324 691 333
rect 717 327 719 339
rect 724 327 726 339
rect 734 327 736 336
rect 744 327 746 336
rect 760 322 762 331
rect 781 324 783 335
rect 788 324 790 335
rect 801 324 803 333
rect 848 324 850 335
rect 855 324 857 335
rect 868 324 870 333
rect 888 324 890 335
rect 895 324 897 335
rect 908 324 910 333
rect 936 327 938 339
rect 943 327 945 339
rect 953 327 955 336
rect 963 327 965 336
rect 979 322 981 331
rect 1000 324 1002 335
rect 1007 324 1009 335
rect 1020 324 1022 333
rect 208 219 210 228
rect 221 217 223 228
rect 228 217 230 228
rect 248 217 250 228
rect 255 217 257 228
rect 268 219 270 228
rect 288 219 290 228
rect 301 217 303 228
rect 308 217 310 228
rect 329 221 331 230
rect 345 216 347 225
rect 355 216 357 225
rect 365 213 367 225
rect 372 213 374 225
rect 424 219 426 228
rect 437 217 439 228
rect 444 217 446 228
rect 464 217 466 228
rect 471 217 473 228
rect 484 219 486 228
rect 504 219 506 228
rect 517 217 519 228
rect 524 217 526 228
rect 545 221 547 230
rect 561 216 563 225
rect 571 216 573 225
rect 581 213 583 225
rect 588 213 590 225
rect 629 219 631 228
rect 642 217 644 228
rect 649 217 651 228
rect 669 217 671 228
rect 676 217 678 228
rect 689 219 691 228
rect 709 219 711 228
rect 722 217 724 228
rect 729 217 731 228
rect 750 221 752 230
rect 766 216 768 225
rect 776 216 778 225
rect 786 213 788 225
rect 793 213 795 225
rect 848 219 850 228
rect 861 217 863 228
rect 868 217 870 228
rect 888 217 890 228
rect 895 217 897 228
rect 908 219 910 228
rect 928 219 930 228
rect 941 217 943 228
rect 948 217 950 228
rect 969 221 971 230
rect 985 216 987 225
rect 995 216 997 225
rect 1005 213 1007 225
rect 1012 213 1014 225
rect 1052 219 1054 228
rect 1065 217 1067 228
rect 1072 217 1074 228
rect 1093 221 1095 230
rect 1109 216 1111 225
rect 1119 216 1121 225
rect 1129 213 1131 225
rect 1136 213 1138 225
rect 158 178 160 187
rect 168 178 170 184
rect 178 178 180 184
rect 198 180 200 189
rect 211 180 213 191
rect 218 180 220 191
rect 239 178 241 187
rect 255 183 257 192
rect 265 183 267 192
rect 275 183 277 195
rect 282 183 284 195
rect 303 180 305 189
rect 316 180 318 191
rect 323 180 325 191
rect 344 178 346 187
rect 360 183 362 192
rect 370 183 372 192
rect 380 183 382 195
rect 387 183 389 195
rect 408 178 410 187
rect 418 178 420 184
rect 428 178 430 184
rect 448 180 450 189
rect 461 180 463 191
rect 468 180 470 191
rect 489 178 491 187
rect 505 183 507 192
rect 515 183 517 192
rect 525 183 527 195
rect 532 183 534 195
rect 553 180 555 189
rect 566 180 568 191
rect 573 180 575 191
rect 594 178 596 187
rect 610 183 612 192
rect 620 183 622 192
rect 630 183 632 195
rect 637 183 639 195
rect 658 178 660 187
rect 668 178 670 184
rect 678 178 680 184
rect 698 180 700 189
rect 711 180 713 191
rect 718 180 720 191
rect 739 178 741 187
rect 755 183 757 192
rect 765 183 767 192
rect 775 183 777 195
rect 782 183 784 195
rect 803 180 805 189
rect 816 180 818 191
rect 823 180 825 191
rect 844 178 846 187
rect 860 183 862 192
rect 870 183 872 192
rect 880 183 882 195
rect 887 183 889 195
rect 908 178 910 187
rect 918 178 920 184
rect 928 178 930 184
rect 948 180 950 189
rect 961 180 963 191
rect 968 180 970 191
rect 989 178 991 187
rect 1005 183 1007 192
rect 1015 183 1017 192
rect 1025 183 1027 195
rect 1032 183 1034 195
rect 1053 180 1055 189
rect 1066 180 1068 191
rect 1073 180 1075 191
rect 1094 178 1096 187
rect 1110 183 1112 192
rect 1120 183 1122 192
rect 1130 183 1132 195
rect 1137 183 1139 195
rect 157 77 159 86
rect 167 80 169 86
rect 177 80 179 86
rect 197 75 199 84
rect 210 73 212 84
rect 217 73 219 84
rect 238 77 240 86
rect 254 72 256 81
rect 264 72 266 81
rect 274 69 276 81
rect 281 69 283 81
rect 302 75 304 84
rect 315 73 317 84
rect 322 73 324 84
rect 343 77 345 86
rect 359 72 361 81
rect 369 72 371 81
rect 379 69 381 81
rect 386 69 388 81
rect 407 77 409 86
rect 417 80 419 86
rect 427 80 429 86
rect 447 75 449 84
rect 460 73 462 84
rect 467 73 469 84
rect 488 77 490 86
rect 504 72 506 81
rect 514 72 516 81
rect 524 69 526 81
rect 531 69 533 81
rect 552 75 554 84
rect 565 73 567 84
rect 572 73 574 84
rect 593 77 595 86
rect 609 72 611 81
rect 619 72 621 81
rect 629 69 631 81
rect 636 69 638 81
rect 657 77 659 86
rect 667 80 669 86
rect 677 80 679 86
rect 697 75 699 84
rect 710 73 712 84
rect 717 73 719 84
rect 738 77 740 86
rect 754 72 756 81
rect 764 72 766 81
rect 774 69 776 81
rect 781 69 783 81
rect 802 75 804 84
rect 815 73 817 84
rect 822 73 824 84
rect 843 77 845 86
rect 859 72 861 81
rect 869 72 871 81
rect 879 69 881 81
rect 886 69 888 81
rect 907 77 909 86
rect 917 80 919 86
rect 927 80 929 86
rect 947 75 949 84
rect 960 73 962 84
rect 967 73 969 84
rect 988 77 990 86
rect 1004 72 1006 81
rect 1014 72 1016 81
rect 1024 69 1026 81
rect 1031 69 1033 81
rect 1052 75 1054 84
rect 1065 73 1067 84
rect 1072 73 1074 84
rect 1093 77 1095 86
rect 1109 72 1111 81
rect 1119 72 1121 81
rect 1129 69 1131 81
rect 1136 69 1138 81
rect 156 34 158 43
rect 166 34 168 40
rect 176 34 178 40
rect 196 36 198 45
rect 209 36 211 47
rect 216 36 218 47
rect 237 34 239 43
rect 253 39 255 48
rect 263 39 265 48
rect 273 39 275 51
rect 280 39 282 51
rect 301 36 303 45
rect 314 36 316 47
rect 321 36 323 47
rect 342 34 344 43
rect 358 39 360 48
rect 368 39 370 48
rect 378 39 380 51
rect 385 39 387 51
rect 406 34 408 43
rect 416 34 418 40
rect 426 34 428 40
rect 446 36 448 45
rect 459 36 461 47
rect 466 36 468 47
rect 487 34 489 43
rect 503 39 505 48
rect 513 39 515 48
rect 523 39 525 51
rect 530 39 532 51
rect 551 36 553 45
rect 564 36 566 47
rect 571 36 573 47
rect 592 34 594 43
rect 608 39 610 48
rect 618 39 620 48
rect 628 39 630 51
rect 635 39 637 51
rect 656 34 658 43
rect 666 34 668 40
rect 676 34 678 40
rect 696 36 698 45
rect 709 36 711 47
rect 716 36 718 47
rect 737 34 739 43
rect 753 39 755 48
rect 763 39 765 48
rect 773 39 775 51
rect 780 39 782 51
rect 801 36 803 45
rect 814 36 816 47
rect 821 36 823 47
rect 842 34 844 43
rect 858 39 860 48
rect 868 39 870 48
rect 878 39 880 51
rect 885 39 887 51
rect 906 34 908 43
rect 916 34 918 40
rect 926 34 928 40
rect 946 36 948 45
rect 959 36 961 47
rect 966 36 968 47
rect 987 34 989 43
rect 1003 39 1005 48
rect 1013 39 1015 48
rect 1023 39 1025 51
rect 1030 39 1032 51
rect 1051 36 1053 45
rect 1064 36 1066 47
rect 1071 36 1073 47
rect 1092 34 1094 43
rect 1108 39 1110 48
rect 1118 39 1120 48
rect 1128 39 1130 51
rect 1135 39 1137 51
<< pmos >>
rect 208 289 210 302
rect 218 289 220 302
rect 228 291 230 309
rect 248 289 250 302
rect 258 289 260 302
rect 268 291 270 309
rect 295 282 297 309
rect 305 291 307 309
rect 315 291 317 309
rect 331 282 333 309
rect 360 289 362 302
rect 370 289 372 302
rect 380 291 382 309
rect 424 289 426 302
rect 434 289 436 302
rect 444 291 446 309
rect 464 289 466 302
rect 474 289 476 302
rect 484 291 486 309
rect 511 282 513 309
rect 521 291 523 309
rect 531 291 533 309
rect 547 282 549 309
rect 576 289 578 302
rect 586 289 588 302
rect 596 291 598 309
rect 629 289 631 302
rect 639 289 641 302
rect 649 291 651 309
rect 669 289 671 302
rect 679 289 681 302
rect 689 291 691 309
rect 716 282 718 309
rect 726 291 728 309
rect 736 291 738 309
rect 752 282 754 309
rect 781 289 783 302
rect 791 289 793 302
rect 801 291 803 309
rect 848 289 850 302
rect 858 289 860 302
rect 868 291 870 309
rect 888 289 890 302
rect 898 289 900 302
rect 908 291 910 309
rect 935 282 937 309
rect 945 291 947 309
rect 955 291 957 309
rect 971 282 973 309
rect 1000 289 1002 302
rect 1010 289 1012 302
rect 1020 291 1022 309
rect 208 243 210 261
rect 218 250 220 263
rect 228 250 230 263
rect 248 250 250 263
rect 258 250 260 263
rect 268 243 270 261
rect 288 243 290 261
rect 298 250 300 263
rect 308 250 310 263
rect 337 243 339 270
rect 353 243 355 261
rect 363 243 365 261
rect 373 243 375 270
rect 424 243 426 261
rect 434 250 436 263
rect 444 250 446 263
rect 464 250 466 263
rect 474 250 476 263
rect 484 243 486 261
rect 504 243 506 261
rect 514 250 516 263
rect 524 250 526 263
rect 553 243 555 270
rect 569 243 571 261
rect 579 243 581 261
rect 589 243 591 270
rect 629 243 631 261
rect 639 250 641 263
rect 649 250 651 263
rect 669 250 671 263
rect 679 250 681 263
rect 689 243 691 261
rect 709 243 711 261
rect 719 250 721 263
rect 729 250 731 263
rect 758 243 760 270
rect 774 243 776 261
rect 784 243 786 261
rect 794 243 796 270
rect 848 243 850 261
rect 858 250 860 263
rect 868 250 870 263
rect 888 250 890 263
rect 898 250 900 263
rect 908 243 910 261
rect 928 243 930 261
rect 938 250 940 263
rect 948 250 950 263
rect 977 243 979 270
rect 993 243 995 261
rect 1003 243 1005 261
rect 1013 243 1015 270
rect 1052 243 1054 261
rect 1062 250 1064 263
rect 1072 250 1074 263
rect 1101 243 1103 270
rect 1117 243 1119 261
rect 1127 243 1129 261
rect 1137 243 1139 270
rect 158 148 160 166
rect 171 138 173 159
rect 178 138 180 159
rect 198 147 200 165
rect 208 145 210 158
rect 218 145 220 158
rect 247 138 249 165
rect 263 147 265 165
rect 273 147 275 165
rect 283 138 285 165
rect 303 147 305 165
rect 313 145 315 158
rect 323 145 325 158
rect 352 138 354 165
rect 368 147 370 165
rect 378 147 380 165
rect 388 138 390 165
rect 408 148 410 166
rect 421 138 423 159
rect 428 138 430 159
rect 448 147 450 165
rect 458 145 460 158
rect 468 145 470 158
rect 497 138 499 165
rect 513 147 515 165
rect 523 147 525 165
rect 533 138 535 165
rect 553 147 555 165
rect 563 145 565 158
rect 573 145 575 158
rect 602 138 604 165
rect 618 147 620 165
rect 628 147 630 165
rect 638 138 640 165
rect 658 148 660 166
rect 671 138 673 159
rect 678 138 680 159
rect 698 147 700 165
rect 708 145 710 158
rect 718 145 720 158
rect 747 138 749 165
rect 763 147 765 165
rect 773 147 775 165
rect 783 138 785 165
rect 803 147 805 165
rect 813 145 815 158
rect 823 145 825 158
rect 852 138 854 165
rect 868 147 870 165
rect 878 147 880 165
rect 888 138 890 165
rect 908 148 910 166
rect 921 138 923 159
rect 928 138 930 159
rect 948 147 950 165
rect 958 145 960 158
rect 968 145 970 158
rect 997 138 999 165
rect 1013 147 1015 165
rect 1023 147 1025 165
rect 1033 138 1035 165
rect 1053 147 1055 165
rect 1063 145 1065 158
rect 1073 145 1075 158
rect 1102 138 1104 165
rect 1118 147 1120 165
rect 1128 147 1130 165
rect 1138 138 1140 165
rect 157 98 159 116
rect 170 105 172 126
rect 177 105 179 126
rect 197 99 199 117
rect 207 106 209 119
rect 217 106 219 119
rect 246 99 248 126
rect 262 99 264 117
rect 272 99 274 117
rect 282 99 284 126
rect 302 99 304 117
rect 312 106 314 119
rect 322 106 324 119
rect 351 99 353 126
rect 367 99 369 117
rect 377 99 379 117
rect 387 99 389 126
rect 407 98 409 116
rect 420 105 422 126
rect 427 105 429 126
rect 447 99 449 117
rect 457 106 459 119
rect 467 106 469 119
rect 496 99 498 126
rect 512 99 514 117
rect 522 99 524 117
rect 532 99 534 126
rect 552 99 554 117
rect 562 106 564 119
rect 572 106 574 119
rect 601 99 603 126
rect 617 99 619 117
rect 627 99 629 117
rect 637 99 639 126
rect 657 98 659 116
rect 670 105 672 126
rect 677 105 679 126
rect 697 99 699 117
rect 707 106 709 119
rect 717 106 719 119
rect 746 99 748 126
rect 762 99 764 117
rect 772 99 774 117
rect 782 99 784 126
rect 802 99 804 117
rect 812 106 814 119
rect 822 106 824 119
rect 851 99 853 126
rect 867 99 869 117
rect 877 99 879 117
rect 887 99 889 126
rect 907 98 909 116
rect 920 105 922 126
rect 927 105 929 126
rect 947 99 949 117
rect 957 106 959 119
rect 967 106 969 119
rect 996 99 998 126
rect 1012 99 1014 117
rect 1022 99 1024 117
rect 1032 99 1034 126
rect 1052 99 1054 117
rect 1062 106 1064 119
rect 1072 106 1074 119
rect 1101 99 1103 126
rect 1117 99 1119 117
rect 1127 99 1129 117
rect 1137 99 1139 126
rect 156 4 158 22
rect 169 -6 171 15
rect 176 -6 178 15
rect 196 3 198 21
rect 206 1 208 14
rect 216 1 218 14
rect 245 -6 247 21
rect 261 3 263 21
rect 271 3 273 21
rect 281 -6 283 21
rect 301 3 303 21
rect 311 1 313 14
rect 321 1 323 14
rect 350 -6 352 21
rect 366 3 368 21
rect 376 3 378 21
rect 386 -6 388 21
rect 406 4 408 22
rect 419 -6 421 15
rect 426 -6 428 15
rect 446 3 448 21
rect 456 1 458 14
rect 466 1 468 14
rect 495 -6 497 21
rect 511 3 513 21
rect 521 3 523 21
rect 531 -6 533 21
rect 551 3 553 21
rect 561 1 563 14
rect 571 1 573 14
rect 600 -6 602 21
rect 616 3 618 21
rect 626 3 628 21
rect 636 -6 638 21
rect 656 4 658 22
rect 669 -6 671 15
rect 676 -6 678 15
rect 696 3 698 21
rect 706 1 708 14
rect 716 1 718 14
rect 745 -6 747 21
rect 761 3 763 21
rect 771 3 773 21
rect 781 -6 783 21
rect 801 3 803 21
rect 811 1 813 14
rect 821 1 823 14
rect 850 -6 852 21
rect 866 3 868 21
rect 876 3 878 21
rect 886 -6 888 21
rect 906 4 908 22
rect 919 -6 921 15
rect 926 -6 928 15
rect 946 3 948 21
rect 956 1 958 14
rect 966 1 968 14
rect 995 -6 997 21
rect 1011 3 1013 21
rect 1021 3 1023 21
rect 1031 -6 1033 21
rect 1051 3 1053 21
rect 1061 1 1063 14
rect 1071 1 1073 14
rect 1100 -6 1102 21
rect 1116 3 1118 21
rect 1126 3 1128 21
rect 1136 -6 1138 21
<< polyct0 >>
rect 226 315 228 317
rect 266 315 268 317
rect 297 314 299 316
rect 307 315 309 317
rect 378 315 380 317
rect 442 315 444 317
rect 482 315 484 317
rect 513 314 515 316
rect 523 315 525 317
rect 594 315 596 317
rect 647 315 649 317
rect 687 315 689 317
rect 718 314 720 316
rect 728 315 730 317
rect 799 315 801 317
rect 866 315 868 317
rect 906 315 908 317
rect 937 314 939 316
rect 947 315 949 317
rect 1018 315 1020 317
rect 210 235 212 237
rect 266 235 268 237
rect 290 235 292 237
rect 361 235 363 237
rect 371 236 373 238
rect 426 235 428 237
rect 482 235 484 237
rect 506 235 508 237
rect 577 235 579 237
rect 587 236 589 238
rect 631 235 633 237
rect 687 235 689 237
rect 711 235 713 237
rect 782 235 784 237
rect 792 236 794 238
rect 850 235 852 237
rect 906 235 908 237
rect 930 235 932 237
rect 1001 235 1003 237
rect 1011 236 1013 238
rect 1054 235 1056 237
rect 1125 235 1127 237
rect 1135 236 1137 238
rect 160 171 162 173
rect 200 171 202 173
rect 271 171 273 173
rect 281 170 283 172
rect 305 171 307 173
rect 376 171 378 173
rect 386 170 388 172
rect 410 171 412 173
rect 450 171 452 173
rect 521 171 523 173
rect 531 170 533 172
rect 555 171 557 173
rect 626 171 628 173
rect 636 170 638 172
rect 660 171 662 173
rect 700 171 702 173
rect 771 171 773 173
rect 781 170 783 172
rect 805 171 807 173
rect 876 171 878 173
rect 886 170 888 172
rect 910 171 912 173
rect 950 171 952 173
rect 1021 171 1023 173
rect 1031 170 1033 172
rect 1055 171 1057 173
rect 1126 171 1128 173
rect 1136 170 1138 172
rect 159 91 161 93
rect 199 91 201 93
rect 270 91 272 93
rect 280 92 282 94
rect 304 91 306 93
rect 375 91 377 93
rect 385 92 387 94
rect 409 91 411 93
rect 449 91 451 93
rect 520 91 522 93
rect 530 92 532 94
rect 554 91 556 93
rect 625 91 627 93
rect 635 92 637 94
rect 659 91 661 93
rect 699 91 701 93
rect 770 91 772 93
rect 780 92 782 94
rect 804 91 806 93
rect 875 91 877 93
rect 885 92 887 94
rect 909 91 911 93
rect 949 91 951 93
rect 1020 91 1022 93
rect 1030 92 1032 94
rect 1054 91 1056 93
rect 1125 91 1127 93
rect 1135 92 1137 94
rect 158 27 160 29
rect 198 27 200 29
rect 269 27 271 29
rect 279 26 281 28
rect 303 27 305 29
rect 374 27 376 29
rect 384 26 386 28
rect 408 27 410 29
rect 448 27 450 29
rect 519 27 521 29
rect 529 26 531 28
rect 553 27 555 29
rect 624 27 626 29
rect 634 26 636 28
rect 658 27 660 29
rect 698 27 700 29
rect 769 27 771 29
rect 779 26 781 28
rect 803 27 805 29
rect 874 27 876 29
rect 884 26 886 28
rect 908 27 910 29
rect 948 27 950 29
rect 1019 27 1021 29
rect 1029 26 1031 28
rect 1053 27 1055 29
rect 1124 27 1126 29
rect 1134 26 1136 28
<< polyct1 >>
rect 216 315 218 317
rect 206 307 208 309
rect 256 315 258 317
rect 328 320 330 322
rect 246 307 248 309
rect 368 315 370 317
rect 344 307 346 309
rect 358 307 360 309
rect 432 315 434 317
rect 422 307 424 309
rect 472 315 474 317
rect 544 320 546 322
rect 462 307 464 309
rect 584 315 586 317
rect 560 307 562 309
rect 574 307 576 309
rect 637 315 639 317
rect 627 307 629 309
rect 677 315 679 317
rect 749 320 751 322
rect 667 307 669 309
rect 789 315 791 317
rect 765 307 767 309
rect 779 307 781 309
rect 856 315 858 317
rect 846 307 848 309
rect 896 315 898 317
rect 968 320 970 322
rect 886 307 888 309
rect 1008 315 1010 317
rect 984 307 986 309
rect 998 307 1000 309
rect 230 243 232 245
rect 246 243 248 245
rect 220 235 222 237
rect 256 235 258 237
rect 310 243 312 245
rect 324 243 326 245
rect 300 235 302 237
rect 446 243 448 245
rect 462 243 464 245
rect 340 230 342 232
rect 436 235 438 237
rect 472 235 474 237
rect 526 243 528 245
rect 540 243 542 245
rect 516 235 518 237
rect 651 243 653 245
rect 667 243 669 245
rect 556 230 558 232
rect 641 235 643 237
rect 677 235 679 237
rect 731 243 733 245
rect 745 243 747 245
rect 721 235 723 237
rect 870 243 872 245
rect 886 243 888 245
rect 761 230 763 232
rect 860 235 862 237
rect 896 235 898 237
rect 950 243 952 245
rect 964 243 966 245
rect 940 235 942 237
rect 1074 243 1076 245
rect 1088 243 1090 245
rect 980 230 982 232
rect 1064 235 1066 237
rect 1104 230 1106 232
rect 170 171 172 173
rect 210 171 212 173
rect 180 164 182 166
rect 250 176 252 178
rect 220 163 222 165
rect 315 171 317 173
rect 234 163 236 165
rect 355 176 357 178
rect 325 163 327 165
rect 420 171 422 173
rect 339 163 341 165
rect 460 171 462 173
rect 430 164 432 166
rect 500 176 502 178
rect 470 163 472 165
rect 565 171 567 173
rect 484 163 486 165
rect 605 176 607 178
rect 575 163 577 165
rect 670 171 672 173
rect 589 163 591 165
rect 710 171 712 173
rect 680 164 682 166
rect 750 176 752 178
rect 720 163 722 165
rect 815 171 817 173
rect 734 163 736 165
rect 855 176 857 178
rect 825 163 827 165
rect 920 171 922 173
rect 839 163 841 165
rect 960 171 962 173
rect 930 164 932 166
rect 1000 176 1002 178
rect 970 163 972 165
rect 1065 171 1067 173
rect 984 163 986 165
rect 1105 176 1107 178
rect 1075 163 1077 165
rect 1089 163 1091 165
rect 179 98 181 100
rect 169 91 171 93
rect 219 99 221 101
rect 233 99 235 101
rect 209 91 211 93
rect 324 99 326 101
rect 338 99 340 101
rect 249 86 251 88
rect 314 91 316 93
rect 429 98 431 100
rect 354 86 356 88
rect 419 91 421 93
rect 469 99 471 101
rect 483 99 485 101
rect 459 91 461 93
rect 574 99 576 101
rect 588 99 590 101
rect 499 86 501 88
rect 564 91 566 93
rect 679 98 681 100
rect 604 86 606 88
rect 669 91 671 93
rect 719 99 721 101
rect 733 99 735 101
rect 709 91 711 93
rect 824 99 826 101
rect 838 99 840 101
rect 749 86 751 88
rect 814 91 816 93
rect 929 98 931 100
rect 854 86 856 88
rect 919 91 921 93
rect 969 99 971 101
rect 983 99 985 101
rect 959 91 961 93
rect 1074 99 1076 101
rect 1088 99 1090 101
rect 999 86 1001 88
rect 1064 91 1066 93
rect 1104 86 1106 88
rect 168 27 170 29
rect 208 27 210 29
rect 178 20 180 22
rect 248 32 250 34
rect 218 19 220 21
rect 313 27 315 29
rect 232 19 234 21
rect 353 32 355 34
rect 323 19 325 21
rect 418 27 420 29
rect 337 19 339 21
rect 458 27 460 29
rect 428 20 430 22
rect 498 32 500 34
rect 468 19 470 21
rect 563 27 565 29
rect 482 19 484 21
rect 603 32 605 34
rect 573 19 575 21
rect 668 27 670 29
rect 587 19 589 21
rect 708 27 710 29
rect 678 20 680 22
rect 748 32 750 34
rect 718 19 720 21
rect 813 27 815 29
rect 732 19 734 21
rect 853 32 855 34
rect 823 19 825 21
rect 918 27 920 29
rect 837 19 839 21
rect 958 27 960 29
rect 928 20 930 22
rect 998 32 1000 34
rect 968 19 970 21
rect 1063 27 1065 29
rect 982 19 984 21
rect 1103 32 1105 34
rect 1073 19 1075 21
rect 1087 19 1089 21
<< ndifct0 >>
rect 203 331 205 333
rect 243 331 245 333
rect 318 329 320 331
rect 330 332 332 334
rect 355 331 357 333
rect 344 324 346 326
rect 419 331 421 333
rect 459 331 461 333
rect 534 329 536 331
rect 546 332 548 334
rect 571 331 573 333
rect 560 324 562 326
rect 624 331 626 333
rect 664 331 666 333
rect 739 329 741 331
rect 751 332 753 334
rect 776 331 778 333
rect 765 324 767 326
rect 843 331 845 333
rect 883 331 885 333
rect 958 329 960 331
rect 970 332 972 334
rect 995 331 997 333
rect 984 324 986 326
rect 233 219 235 221
rect 243 219 245 221
rect 324 226 326 228
rect 313 219 315 221
rect 338 218 340 220
rect 350 221 352 223
rect 449 219 451 221
rect 459 219 461 221
rect 540 226 542 228
rect 529 219 531 221
rect 554 218 556 220
rect 566 221 568 223
rect 654 219 656 221
rect 664 219 666 221
rect 745 226 747 228
rect 734 219 736 221
rect 759 218 761 220
rect 771 221 773 223
rect 873 219 875 221
rect 883 219 885 221
rect 964 226 966 228
rect 953 219 955 221
rect 978 218 980 220
rect 990 221 992 223
rect 1088 226 1090 228
rect 1077 219 1079 221
rect 1102 218 1104 220
rect 1114 221 1116 223
rect 164 193 166 195
rect 183 193 185 195
rect 173 180 175 182
rect 223 187 225 189
rect 248 188 250 190
rect 234 180 236 182
rect 260 185 262 187
rect 328 187 330 189
rect 353 188 355 190
rect 339 180 341 182
rect 365 185 367 187
rect 414 193 416 195
rect 433 193 435 195
rect 423 180 425 182
rect 473 187 475 189
rect 498 188 500 190
rect 484 180 486 182
rect 510 185 512 187
rect 578 187 580 189
rect 603 188 605 190
rect 589 180 591 182
rect 615 185 617 187
rect 664 193 666 195
rect 683 193 685 195
rect 673 180 675 182
rect 723 187 725 189
rect 748 188 750 190
rect 734 180 736 182
rect 760 185 762 187
rect 828 187 830 189
rect 853 188 855 190
rect 839 180 841 182
rect 865 185 867 187
rect 914 193 916 195
rect 933 193 935 195
rect 923 180 925 182
rect 973 187 975 189
rect 998 188 1000 190
rect 984 180 986 182
rect 1010 185 1012 187
rect 1078 187 1080 189
rect 1103 188 1105 190
rect 1089 180 1091 182
rect 1115 185 1117 187
rect 172 82 174 84
rect 163 69 165 71
rect 233 82 235 84
rect 222 75 224 77
rect 247 74 249 76
rect 182 69 184 71
rect 259 77 261 79
rect 338 82 340 84
rect 327 75 329 77
rect 352 74 354 76
rect 364 77 366 79
rect 422 82 424 84
rect 413 69 415 71
rect 483 82 485 84
rect 472 75 474 77
rect 497 74 499 76
rect 432 69 434 71
rect 509 77 511 79
rect 588 82 590 84
rect 577 75 579 77
rect 602 74 604 76
rect 614 77 616 79
rect 672 82 674 84
rect 663 69 665 71
rect 733 82 735 84
rect 722 75 724 77
rect 747 74 749 76
rect 682 69 684 71
rect 759 77 761 79
rect 838 82 840 84
rect 827 75 829 77
rect 852 74 854 76
rect 864 77 866 79
rect 922 82 924 84
rect 913 69 915 71
rect 983 82 985 84
rect 972 75 974 77
rect 997 74 999 76
rect 932 69 934 71
rect 1009 77 1011 79
rect 1088 82 1090 84
rect 1077 75 1079 77
rect 1102 74 1104 76
rect 1114 77 1116 79
rect 162 49 164 51
rect 181 49 183 51
rect 171 36 173 38
rect 221 43 223 45
rect 246 44 248 46
rect 232 36 234 38
rect 258 41 260 43
rect 326 43 328 45
rect 351 44 353 46
rect 337 36 339 38
rect 363 41 365 43
rect 412 49 414 51
rect 431 49 433 51
rect 421 36 423 38
rect 471 43 473 45
rect 496 44 498 46
rect 482 36 484 38
rect 508 41 510 43
rect 576 43 578 45
rect 601 44 603 46
rect 587 36 589 38
rect 613 41 615 43
rect 662 49 664 51
rect 681 49 683 51
rect 671 36 673 38
rect 721 43 723 45
rect 746 44 748 46
rect 732 36 734 38
rect 758 41 760 43
rect 826 43 828 45
rect 851 44 853 46
rect 837 36 839 38
rect 863 41 865 43
rect 912 49 914 51
rect 931 49 933 51
rect 921 36 923 38
rect 971 43 973 45
rect 996 44 998 46
rect 982 36 984 38
rect 1008 41 1010 43
rect 1076 43 1078 45
rect 1101 44 1103 46
rect 1087 36 1089 38
rect 1113 41 1115 43
<< ndifct1 >>
rect 222 341 224 343
rect 262 341 264 343
rect 290 341 292 343
rect 233 329 235 331
rect 273 329 275 331
rect 374 341 376 343
rect 308 331 310 333
rect 438 341 440 343
rect 478 341 480 343
rect 385 329 387 331
rect 506 341 508 343
rect 449 329 451 331
rect 489 329 491 331
rect 590 341 592 343
rect 524 331 526 333
rect 643 341 645 343
rect 683 341 685 343
rect 601 329 603 331
rect 711 341 713 343
rect 654 329 656 331
rect 694 329 696 331
rect 795 341 797 343
rect 729 331 731 333
rect 862 341 864 343
rect 902 341 904 343
rect 806 329 808 331
rect 930 341 932 343
rect 873 329 875 331
rect 913 329 915 331
rect 1014 341 1016 343
rect 948 331 950 333
rect 1025 329 1027 331
rect 203 221 205 223
rect 273 221 275 223
rect 283 221 285 223
rect 214 209 216 211
rect 262 209 264 211
rect 360 219 362 221
rect 294 209 296 211
rect 419 221 421 223
rect 489 221 491 223
rect 499 221 501 223
rect 378 209 380 211
rect 430 209 432 211
rect 478 209 480 211
rect 576 219 578 221
rect 510 209 512 211
rect 624 221 626 223
rect 694 221 696 223
rect 704 221 706 223
rect 594 209 596 211
rect 635 209 637 211
rect 683 209 685 211
rect 781 219 783 221
rect 715 209 717 211
rect 843 221 845 223
rect 913 221 915 223
rect 923 221 925 223
rect 799 209 801 211
rect 854 209 856 211
rect 902 209 904 211
rect 1000 219 1002 221
rect 934 209 936 211
rect 1047 221 1049 223
rect 1018 209 1020 211
rect 1124 219 1126 221
rect 1058 209 1060 211
rect 1142 209 1144 211
rect 204 197 206 199
rect 153 180 155 182
rect 288 197 290 199
rect 309 197 311 199
rect 193 185 195 187
rect 270 187 272 189
rect 393 197 395 199
rect 298 185 300 187
rect 375 187 377 189
rect 454 197 456 199
rect 403 180 405 182
rect 538 197 540 199
rect 559 197 561 199
rect 443 185 445 187
rect 520 187 522 189
rect 643 197 645 199
rect 548 185 550 187
rect 625 187 627 189
rect 704 197 706 199
rect 653 180 655 182
rect 788 197 790 199
rect 809 197 811 199
rect 693 185 695 187
rect 770 187 772 189
rect 893 197 895 199
rect 798 185 800 187
rect 875 187 877 189
rect 954 197 956 199
rect 903 180 905 182
rect 1038 197 1040 199
rect 1059 197 1061 199
rect 943 185 945 187
rect 1020 187 1022 189
rect 1143 197 1145 199
rect 1048 185 1050 187
rect 1125 187 1127 189
rect 152 82 154 84
rect 192 77 194 79
rect 269 75 271 77
rect 203 65 205 67
rect 297 77 299 79
rect 402 82 404 84
rect 287 65 289 67
rect 374 75 376 77
rect 308 65 310 67
rect 442 77 444 79
rect 392 65 394 67
rect 519 75 521 77
rect 453 65 455 67
rect 547 77 549 79
rect 652 82 654 84
rect 537 65 539 67
rect 624 75 626 77
rect 558 65 560 67
rect 692 77 694 79
rect 642 65 644 67
rect 769 75 771 77
rect 703 65 705 67
rect 797 77 799 79
rect 902 82 904 84
rect 787 65 789 67
rect 874 75 876 77
rect 808 65 810 67
rect 942 77 944 79
rect 892 65 894 67
rect 1019 75 1021 77
rect 953 65 955 67
rect 1047 77 1049 79
rect 1037 65 1039 67
rect 1124 75 1126 77
rect 1058 65 1060 67
rect 1142 65 1144 67
rect 202 53 204 55
rect 151 36 153 38
rect 286 53 288 55
rect 307 53 309 55
rect 191 41 193 43
rect 268 43 270 45
rect 391 53 393 55
rect 296 41 298 43
rect 373 43 375 45
rect 452 53 454 55
rect 401 36 403 38
rect 536 53 538 55
rect 557 53 559 55
rect 441 41 443 43
rect 518 43 520 45
rect 641 53 643 55
rect 546 41 548 43
rect 623 43 625 45
rect 702 53 704 55
rect 651 36 653 38
rect 786 53 788 55
rect 807 53 809 55
rect 691 41 693 43
rect 768 43 770 45
rect 891 53 893 55
rect 796 41 798 43
rect 873 43 875 45
rect 952 53 954 55
rect 901 36 903 38
rect 1036 53 1038 55
rect 1057 53 1059 55
rect 941 41 943 43
rect 1018 43 1020 45
rect 1141 53 1143 55
rect 1046 41 1048 43
rect 1123 43 1125 45
<< ntiect1 >>
rect 232 281 234 283
rect 272 281 274 283
rect 310 281 312 283
rect 384 281 386 283
rect 448 281 450 283
rect 488 281 490 283
rect 526 281 528 283
rect 600 281 602 283
rect 653 281 655 283
rect 693 281 695 283
rect 731 281 733 283
rect 805 281 807 283
rect 872 281 874 283
rect 912 281 914 283
rect 950 281 952 283
rect 1024 281 1026 283
rect 204 269 206 271
rect 272 269 274 271
rect 284 269 286 271
rect 358 269 360 271
rect 420 269 422 271
rect 488 269 490 271
rect 500 269 502 271
rect 574 269 576 271
rect 625 269 627 271
rect 693 269 695 271
rect 705 269 707 271
rect 779 269 781 271
rect 844 269 846 271
rect 912 269 914 271
rect 924 269 926 271
rect 998 269 1000 271
rect 1048 269 1050 271
rect 1122 269 1124 271
rect 154 137 156 139
rect 194 137 196 139
rect 268 137 270 139
rect 299 137 301 139
rect 373 137 375 139
rect 404 137 406 139
rect 444 137 446 139
rect 518 137 520 139
rect 549 137 551 139
rect 623 137 625 139
rect 654 137 656 139
rect 694 137 696 139
rect 768 137 770 139
rect 799 137 801 139
rect 873 137 875 139
rect 904 137 906 139
rect 944 137 946 139
rect 1018 137 1020 139
rect 1049 137 1051 139
rect 1123 137 1125 139
rect 153 125 155 127
rect 193 125 195 127
rect 267 125 269 127
rect 298 125 300 127
rect 372 125 374 127
rect 403 125 405 127
rect 443 125 445 127
rect 517 125 519 127
rect 548 125 550 127
rect 622 125 624 127
rect 653 125 655 127
rect 693 125 695 127
rect 767 125 769 127
rect 798 125 800 127
rect 872 125 874 127
rect 903 125 905 127
rect 943 125 945 127
rect 1017 125 1019 127
rect 1048 125 1050 127
rect 1122 125 1124 127
rect 152 -7 154 -5
rect 192 -7 194 -5
rect 266 -7 268 -5
rect 297 -7 299 -5
rect 371 -7 373 -5
rect 402 -7 404 -5
rect 442 -7 444 -5
rect 516 -7 518 -5
rect 547 -7 549 -5
rect 621 -7 623 -5
rect 652 -7 654 -5
rect 692 -7 694 -5
rect 766 -7 768 -5
rect 797 -7 799 -5
rect 871 -7 873 -5
rect 902 -7 904 -5
rect 942 -7 944 -5
rect 1016 -7 1018 -5
rect 1047 -7 1049 -5
rect 1121 -7 1123 -5
<< ptiect1 >>
rect 232 341 234 343
rect 272 341 274 343
rect 343 341 345 343
rect 384 341 386 343
rect 448 341 450 343
rect 488 341 490 343
rect 559 341 561 343
rect 600 341 602 343
rect 653 341 655 343
rect 693 341 695 343
rect 764 341 766 343
rect 805 341 807 343
rect 872 341 874 343
rect 912 341 914 343
rect 983 341 985 343
rect 1024 341 1026 343
rect 204 209 206 211
rect 272 209 274 211
rect 284 209 286 211
rect 325 209 327 211
rect 420 209 422 211
rect 488 209 490 211
rect 500 209 502 211
rect 541 209 543 211
rect 625 209 627 211
rect 693 209 695 211
rect 705 209 707 211
rect 746 209 748 211
rect 844 209 846 211
rect 912 209 914 211
rect 924 209 926 211
rect 965 209 967 211
rect 1048 209 1050 211
rect 1089 209 1091 211
rect 154 197 156 199
rect 194 197 196 199
rect 235 197 237 199
rect 299 197 301 199
rect 340 197 342 199
rect 404 197 406 199
rect 444 197 446 199
rect 485 197 487 199
rect 549 197 551 199
rect 590 197 592 199
rect 654 197 656 199
rect 694 197 696 199
rect 735 197 737 199
rect 799 197 801 199
rect 840 197 842 199
rect 904 197 906 199
rect 944 197 946 199
rect 985 197 987 199
rect 1049 197 1051 199
rect 1090 197 1092 199
rect 153 65 155 67
rect 193 65 195 67
rect 234 65 236 67
rect 298 65 300 67
rect 339 65 341 67
rect 403 65 405 67
rect 443 65 445 67
rect 484 65 486 67
rect 548 65 550 67
rect 589 65 591 67
rect 653 65 655 67
rect 693 65 695 67
rect 734 65 736 67
rect 798 65 800 67
rect 839 65 841 67
rect 903 65 905 67
rect 943 65 945 67
rect 984 65 986 67
rect 1048 65 1050 67
rect 1089 65 1091 67
rect 152 53 154 55
rect 192 53 194 55
rect 233 53 235 55
rect 297 53 299 55
rect 338 53 340 55
rect 402 53 404 55
rect 442 53 444 55
rect 483 53 485 55
rect 547 53 549 55
rect 588 53 590 55
rect 652 53 654 55
rect 692 53 694 55
rect 733 53 735 55
rect 797 53 799 55
rect 838 53 840 55
rect 902 53 904 55
rect 942 53 944 55
rect 983 53 985 55
rect 1047 53 1049 55
rect 1088 53 1090 55
<< pdifct0 >>
rect 203 291 205 293
rect 213 298 215 300
rect 213 291 215 293
rect 223 293 225 295
rect 243 291 245 293
rect 253 298 255 300
rect 253 291 255 293
rect 263 293 265 295
rect 290 290 292 292
rect 310 305 312 307
rect 310 298 312 300
rect 326 291 328 293
rect 326 284 328 286
rect 336 305 338 307
rect 355 291 357 293
rect 365 298 367 300
rect 365 291 367 293
rect 375 293 377 295
rect 419 291 421 293
rect 429 298 431 300
rect 429 291 431 293
rect 439 293 441 295
rect 459 291 461 293
rect 469 298 471 300
rect 469 291 471 293
rect 479 293 481 295
rect 506 290 508 292
rect 526 305 528 307
rect 526 298 528 300
rect 542 291 544 293
rect 542 284 544 286
rect 552 305 554 307
rect 571 291 573 293
rect 581 298 583 300
rect 581 291 583 293
rect 591 293 593 295
rect 624 291 626 293
rect 634 298 636 300
rect 634 291 636 293
rect 644 293 646 295
rect 664 291 666 293
rect 674 298 676 300
rect 674 291 676 293
rect 684 293 686 295
rect 711 290 713 292
rect 731 305 733 307
rect 731 298 733 300
rect 747 291 749 293
rect 747 284 749 286
rect 757 305 759 307
rect 776 291 778 293
rect 786 298 788 300
rect 786 291 788 293
rect 796 293 798 295
rect 843 291 845 293
rect 853 298 855 300
rect 853 291 855 293
rect 863 293 865 295
rect 883 291 885 293
rect 893 298 895 300
rect 893 291 895 293
rect 903 293 905 295
rect 930 290 932 292
rect 950 305 952 307
rect 950 298 952 300
rect 966 291 968 293
rect 966 284 968 286
rect 976 305 978 307
rect 995 291 997 293
rect 1005 298 1007 300
rect 1005 291 1007 293
rect 1015 293 1017 295
rect 213 257 215 259
rect 223 259 225 261
rect 223 252 225 254
rect 233 259 235 261
rect 243 259 245 261
rect 253 259 255 261
rect 253 252 255 254
rect 263 257 265 259
rect 293 257 295 259
rect 303 259 305 261
rect 303 252 305 254
rect 313 259 315 261
rect 332 245 334 247
rect 342 266 344 268
rect 342 259 344 261
rect 358 252 360 254
rect 358 245 360 247
rect 378 260 380 262
rect 429 257 431 259
rect 439 259 441 261
rect 439 252 441 254
rect 449 259 451 261
rect 459 259 461 261
rect 469 259 471 261
rect 469 252 471 254
rect 479 257 481 259
rect 509 257 511 259
rect 519 259 521 261
rect 519 252 521 254
rect 529 259 531 261
rect 548 245 550 247
rect 558 266 560 268
rect 558 259 560 261
rect 574 252 576 254
rect 574 245 576 247
rect 594 260 596 262
rect 634 257 636 259
rect 644 259 646 261
rect 644 252 646 254
rect 654 259 656 261
rect 664 259 666 261
rect 674 259 676 261
rect 674 252 676 254
rect 684 257 686 259
rect 714 257 716 259
rect 724 259 726 261
rect 724 252 726 254
rect 734 259 736 261
rect 753 245 755 247
rect 763 266 765 268
rect 763 259 765 261
rect 779 252 781 254
rect 779 245 781 247
rect 799 260 801 262
rect 853 257 855 259
rect 863 259 865 261
rect 863 252 865 254
rect 873 259 875 261
rect 883 259 885 261
rect 893 259 895 261
rect 893 252 895 254
rect 903 257 905 259
rect 933 257 935 259
rect 943 259 945 261
rect 943 252 945 254
rect 953 259 955 261
rect 972 245 974 247
rect 982 266 984 268
rect 982 259 984 261
rect 998 252 1000 254
rect 998 245 1000 247
rect 1018 260 1020 262
rect 1057 257 1059 259
rect 1067 259 1069 261
rect 1067 252 1069 254
rect 1077 259 1079 261
rect 1096 245 1098 247
rect 1106 266 1108 268
rect 1106 259 1108 261
rect 1122 252 1124 254
rect 1122 245 1124 247
rect 1142 260 1144 262
rect 164 140 166 142
rect 183 147 185 149
rect 242 161 244 163
rect 203 149 205 151
rect 213 154 215 156
rect 213 147 215 149
rect 223 147 225 149
rect 252 147 254 149
rect 268 161 270 163
rect 268 154 270 156
rect 252 140 254 142
rect 288 146 290 148
rect 347 161 349 163
rect 308 149 310 151
rect 318 154 320 156
rect 318 147 320 149
rect 328 147 330 149
rect 357 147 359 149
rect 373 161 375 163
rect 373 154 375 156
rect 357 140 359 142
rect 393 146 395 148
rect 414 140 416 142
rect 433 147 435 149
rect 492 161 494 163
rect 453 149 455 151
rect 463 154 465 156
rect 463 147 465 149
rect 473 147 475 149
rect 502 147 504 149
rect 518 161 520 163
rect 518 154 520 156
rect 502 140 504 142
rect 538 146 540 148
rect 597 161 599 163
rect 558 149 560 151
rect 568 154 570 156
rect 568 147 570 149
rect 578 147 580 149
rect 607 147 609 149
rect 623 161 625 163
rect 623 154 625 156
rect 607 140 609 142
rect 643 146 645 148
rect 664 140 666 142
rect 683 147 685 149
rect 742 161 744 163
rect 703 149 705 151
rect 713 154 715 156
rect 713 147 715 149
rect 723 147 725 149
rect 752 147 754 149
rect 768 161 770 163
rect 768 154 770 156
rect 752 140 754 142
rect 788 146 790 148
rect 847 161 849 163
rect 808 149 810 151
rect 818 154 820 156
rect 818 147 820 149
rect 828 147 830 149
rect 857 147 859 149
rect 873 161 875 163
rect 873 154 875 156
rect 857 140 859 142
rect 893 146 895 148
rect 914 140 916 142
rect 933 147 935 149
rect 992 161 994 163
rect 953 149 955 151
rect 963 154 965 156
rect 963 147 965 149
rect 973 147 975 149
rect 1002 147 1004 149
rect 1018 161 1020 163
rect 1018 154 1020 156
rect 1002 140 1004 142
rect 1038 146 1040 148
rect 1097 161 1099 163
rect 1058 149 1060 151
rect 1068 154 1070 156
rect 1068 147 1070 149
rect 1078 147 1080 149
rect 1107 147 1109 149
rect 1123 161 1125 163
rect 1123 154 1125 156
rect 1107 140 1109 142
rect 1143 146 1145 148
rect 163 122 165 124
rect 182 115 184 117
rect 202 113 204 115
rect 212 115 214 117
rect 212 108 214 110
rect 222 115 224 117
rect 241 101 243 103
rect 251 122 253 124
rect 251 115 253 117
rect 267 108 269 110
rect 267 101 269 103
rect 287 116 289 118
rect 307 113 309 115
rect 317 115 319 117
rect 317 108 319 110
rect 327 115 329 117
rect 346 101 348 103
rect 356 122 358 124
rect 356 115 358 117
rect 372 108 374 110
rect 372 101 374 103
rect 413 122 415 124
rect 392 116 394 118
rect 432 115 434 117
rect 452 113 454 115
rect 462 115 464 117
rect 462 108 464 110
rect 472 115 474 117
rect 491 101 493 103
rect 501 122 503 124
rect 501 115 503 117
rect 517 108 519 110
rect 517 101 519 103
rect 537 116 539 118
rect 557 113 559 115
rect 567 115 569 117
rect 567 108 569 110
rect 577 115 579 117
rect 596 101 598 103
rect 606 122 608 124
rect 606 115 608 117
rect 622 108 624 110
rect 622 101 624 103
rect 663 122 665 124
rect 642 116 644 118
rect 682 115 684 117
rect 702 113 704 115
rect 712 115 714 117
rect 712 108 714 110
rect 722 115 724 117
rect 741 101 743 103
rect 751 122 753 124
rect 751 115 753 117
rect 767 108 769 110
rect 767 101 769 103
rect 787 116 789 118
rect 807 113 809 115
rect 817 115 819 117
rect 817 108 819 110
rect 827 115 829 117
rect 846 101 848 103
rect 856 122 858 124
rect 856 115 858 117
rect 872 108 874 110
rect 872 101 874 103
rect 913 122 915 124
rect 892 116 894 118
rect 932 115 934 117
rect 952 113 954 115
rect 962 115 964 117
rect 962 108 964 110
rect 972 115 974 117
rect 991 101 993 103
rect 1001 122 1003 124
rect 1001 115 1003 117
rect 1017 108 1019 110
rect 1017 101 1019 103
rect 1037 116 1039 118
rect 1057 113 1059 115
rect 1067 115 1069 117
rect 1067 108 1069 110
rect 1077 115 1079 117
rect 1096 101 1098 103
rect 1106 122 1108 124
rect 1106 115 1108 117
rect 1122 108 1124 110
rect 1122 101 1124 103
rect 1142 116 1144 118
rect 162 -4 164 -2
rect 181 3 183 5
rect 240 17 242 19
rect 201 5 203 7
rect 211 10 213 12
rect 211 3 213 5
rect 221 3 223 5
rect 250 3 252 5
rect 266 17 268 19
rect 266 10 268 12
rect 250 -4 252 -2
rect 286 2 288 4
rect 345 17 347 19
rect 306 5 308 7
rect 316 10 318 12
rect 316 3 318 5
rect 326 3 328 5
rect 355 3 357 5
rect 371 17 373 19
rect 371 10 373 12
rect 355 -4 357 -2
rect 391 2 393 4
rect 412 -4 414 -2
rect 431 3 433 5
rect 490 17 492 19
rect 451 5 453 7
rect 461 10 463 12
rect 461 3 463 5
rect 471 3 473 5
rect 500 3 502 5
rect 516 17 518 19
rect 516 10 518 12
rect 500 -4 502 -2
rect 536 2 538 4
rect 595 17 597 19
rect 556 5 558 7
rect 566 10 568 12
rect 566 3 568 5
rect 576 3 578 5
rect 605 3 607 5
rect 621 17 623 19
rect 621 10 623 12
rect 605 -4 607 -2
rect 641 2 643 4
rect 662 -4 664 -2
rect 681 3 683 5
rect 740 17 742 19
rect 701 5 703 7
rect 711 10 713 12
rect 711 3 713 5
rect 721 3 723 5
rect 750 3 752 5
rect 766 17 768 19
rect 766 10 768 12
rect 750 -4 752 -2
rect 786 2 788 4
rect 845 17 847 19
rect 806 5 808 7
rect 816 10 818 12
rect 816 3 818 5
rect 826 3 828 5
rect 855 3 857 5
rect 871 17 873 19
rect 871 10 873 12
rect 855 -4 857 -2
rect 891 2 893 4
rect 912 -4 914 -2
rect 931 3 933 5
rect 990 17 992 19
rect 951 5 953 7
rect 961 10 963 12
rect 961 3 963 5
rect 971 3 973 5
rect 1000 3 1002 5
rect 1016 17 1018 19
rect 1016 10 1018 12
rect 1000 -4 1002 -2
rect 1036 2 1038 4
rect 1095 17 1097 19
rect 1056 5 1058 7
rect 1066 10 1068 12
rect 1066 3 1068 5
rect 1076 3 1078 5
rect 1105 3 1107 5
rect 1121 17 1123 19
rect 1121 10 1123 12
rect 1105 -4 1107 -2
rect 1141 2 1143 4
<< pdifct1 >>
rect 233 305 235 307
rect 233 298 235 300
rect 273 305 275 307
rect 273 298 275 300
rect 300 298 302 300
rect 385 305 387 307
rect 385 298 387 300
rect 449 305 451 307
rect 449 298 451 300
rect 489 305 491 307
rect 489 298 491 300
rect 516 298 518 300
rect 601 305 603 307
rect 601 298 603 300
rect 654 305 656 307
rect 654 298 656 300
rect 694 305 696 307
rect 694 298 696 300
rect 721 298 723 300
rect 806 305 808 307
rect 806 298 808 300
rect 873 305 875 307
rect 873 298 875 300
rect 913 305 915 307
rect 913 298 915 300
rect 940 298 942 300
rect 1025 305 1027 307
rect 1025 298 1027 300
rect 203 252 205 254
rect 203 245 205 247
rect 273 252 275 254
rect 273 245 275 247
rect 283 252 285 254
rect 283 245 285 247
rect 368 252 370 254
rect 419 252 421 254
rect 419 245 421 247
rect 489 252 491 254
rect 489 245 491 247
rect 499 252 501 254
rect 499 245 501 247
rect 584 252 586 254
rect 624 252 626 254
rect 624 245 626 247
rect 694 252 696 254
rect 694 245 696 247
rect 704 252 706 254
rect 704 245 706 247
rect 789 252 791 254
rect 843 252 845 254
rect 843 245 845 247
rect 913 252 915 254
rect 913 245 915 247
rect 923 252 925 254
rect 923 245 925 247
rect 1008 252 1010 254
rect 1047 252 1049 254
rect 1047 245 1049 247
rect 1132 252 1134 254
rect 153 157 155 159
rect 153 150 155 152
rect 193 161 195 163
rect 193 154 195 156
rect 278 154 280 156
rect 298 161 300 163
rect 298 154 300 156
rect 383 154 385 156
rect 403 157 405 159
rect 403 150 405 152
rect 443 161 445 163
rect 443 154 445 156
rect 528 154 530 156
rect 548 161 550 163
rect 548 154 550 156
rect 633 154 635 156
rect 653 157 655 159
rect 653 150 655 152
rect 693 161 695 163
rect 693 154 695 156
rect 778 154 780 156
rect 798 161 800 163
rect 798 154 800 156
rect 883 154 885 156
rect 903 157 905 159
rect 903 150 905 152
rect 943 161 945 163
rect 943 154 945 156
rect 1028 154 1030 156
rect 1048 161 1050 163
rect 1048 154 1050 156
rect 1133 154 1135 156
rect 152 112 154 114
rect 152 105 154 107
rect 192 108 194 110
rect 192 101 194 103
rect 277 108 279 110
rect 297 108 299 110
rect 297 101 299 103
rect 382 108 384 110
rect 402 112 404 114
rect 402 105 404 107
rect 442 108 444 110
rect 442 101 444 103
rect 527 108 529 110
rect 547 108 549 110
rect 547 101 549 103
rect 632 108 634 110
rect 652 112 654 114
rect 652 105 654 107
rect 692 108 694 110
rect 692 101 694 103
rect 777 108 779 110
rect 797 108 799 110
rect 797 101 799 103
rect 882 108 884 110
rect 902 112 904 114
rect 902 105 904 107
rect 942 108 944 110
rect 942 101 944 103
rect 1027 108 1029 110
rect 1047 108 1049 110
rect 1047 101 1049 103
rect 1132 108 1134 110
rect 151 13 153 15
rect 151 6 153 8
rect 191 17 193 19
rect 191 10 193 12
rect 276 10 278 12
rect 296 17 298 19
rect 296 10 298 12
rect 381 10 383 12
rect 401 13 403 15
rect 401 6 403 8
rect 441 17 443 19
rect 441 10 443 12
rect 526 10 528 12
rect 546 17 548 19
rect 546 10 548 12
rect 631 10 633 12
rect 651 13 653 15
rect 651 6 653 8
rect 691 17 693 19
rect 691 10 693 12
rect 776 10 778 12
rect 796 17 798 19
rect 796 10 798 12
rect 881 10 883 12
rect 901 13 903 15
rect 901 6 903 8
rect 941 17 943 19
rect 941 10 943 12
rect 1026 10 1028 12
rect 1046 17 1048 19
rect 1046 10 1048 12
rect 1131 10 1133 12
<< alu0 >>
rect 201 333 221 334
rect 201 331 203 333
rect 205 331 221 333
rect 201 330 221 331
rect 217 326 221 330
rect 241 333 261 334
rect 241 331 243 333
rect 245 331 261 333
rect 241 330 261 331
rect 232 327 233 329
rect 217 322 229 326
rect 225 317 229 322
rect 225 315 226 317
rect 228 315 229 317
rect 225 303 229 315
rect 257 326 261 330
rect 328 334 334 340
rect 272 327 273 329
rect 257 322 269 326
rect 265 317 269 322
rect 265 315 266 317
rect 268 315 269 317
rect 212 300 229 303
rect 212 298 213 300
rect 215 299 229 300
rect 215 298 216 299
rect 201 293 207 294
rect 201 291 203 293
rect 205 291 207 293
rect 201 284 207 291
rect 212 293 216 298
rect 265 303 269 315
rect 252 300 269 303
rect 252 298 253 300
rect 255 299 269 300
rect 255 298 256 299
rect 212 291 213 293
rect 215 291 216 293
rect 212 289 216 291
rect 221 295 227 296
rect 221 293 223 295
rect 225 293 227 295
rect 221 284 227 293
rect 241 293 247 294
rect 241 291 243 293
rect 245 291 247 293
rect 241 284 247 291
rect 252 293 256 298
rect 317 331 321 333
rect 328 332 330 334
rect 332 332 334 334
rect 328 331 334 332
rect 353 333 373 334
rect 353 331 355 333
rect 357 331 373 333
rect 317 329 318 331
rect 320 329 321 331
rect 353 330 373 331
rect 317 326 321 329
rect 297 322 321 326
rect 297 318 301 322
rect 343 326 347 328
rect 343 324 344 326
rect 346 324 347 326
rect 296 316 301 318
rect 296 314 297 316
rect 299 314 301 316
rect 305 317 321 318
rect 305 315 307 317
rect 309 315 321 317
rect 305 314 321 315
rect 296 312 301 314
rect 297 310 301 312
rect 297 307 313 310
rect 297 306 310 307
rect 309 305 310 306
rect 312 305 313 307
rect 309 300 313 305
rect 309 298 310 300
rect 312 298 313 300
rect 309 296 313 298
rect 317 308 321 314
rect 343 318 347 324
rect 336 314 347 318
rect 369 326 373 330
rect 417 333 437 334
rect 417 331 419 333
rect 421 331 437 333
rect 417 330 437 331
rect 384 327 385 329
rect 369 322 381 326
rect 377 317 381 322
rect 377 315 378 317
rect 380 315 381 317
rect 336 308 340 314
rect 317 307 340 308
rect 317 305 336 307
rect 338 305 340 307
rect 317 304 340 305
rect 252 291 253 293
rect 255 291 256 293
rect 252 289 256 291
rect 261 295 267 296
rect 261 293 263 295
rect 265 293 267 295
rect 317 293 321 304
rect 377 303 381 315
rect 433 326 437 330
rect 457 333 477 334
rect 457 331 459 333
rect 461 331 477 333
rect 457 330 477 331
rect 448 327 449 329
rect 433 322 445 326
rect 441 317 445 322
rect 441 315 442 317
rect 444 315 445 317
rect 364 300 381 303
rect 364 298 365 300
rect 367 299 381 300
rect 367 298 368 299
rect 261 284 267 293
rect 288 292 321 293
rect 288 290 290 292
rect 292 290 321 292
rect 288 289 321 290
rect 325 293 329 295
rect 325 291 326 293
rect 328 291 329 293
rect 325 286 329 291
rect 353 293 359 294
rect 353 291 355 293
rect 357 291 359 293
rect 325 284 326 286
rect 328 284 329 286
rect 353 284 359 291
rect 364 293 368 298
rect 441 303 445 315
rect 473 326 477 330
rect 544 334 550 340
rect 488 327 489 329
rect 473 322 485 326
rect 481 317 485 322
rect 481 315 482 317
rect 484 315 485 317
rect 428 300 445 303
rect 428 298 429 300
rect 431 299 445 300
rect 431 298 432 299
rect 364 291 365 293
rect 367 291 368 293
rect 364 289 368 291
rect 373 295 379 296
rect 373 293 375 295
rect 377 293 379 295
rect 373 284 379 293
rect 417 293 423 294
rect 417 291 419 293
rect 421 291 423 293
rect 417 284 423 291
rect 428 293 432 298
rect 481 303 485 315
rect 468 300 485 303
rect 468 298 469 300
rect 471 299 485 300
rect 471 298 472 299
rect 428 291 429 293
rect 431 291 432 293
rect 428 289 432 291
rect 437 295 443 296
rect 437 293 439 295
rect 441 293 443 295
rect 437 284 443 293
rect 457 293 463 294
rect 457 291 459 293
rect 461 291 463 293
rect 457 284 463 291
rect 468 293 472 298
rect 533 331 537 333
rect 544 332 546 334
rect 548 332 550 334
rect 544 331 550 332
rect 569 333 589 334
rect 569 331 571 333
rect 573 331 589 333
rect 533 329 534 331
rect 536 329 537 331
rect 569 330 589 331
rect 533 326 537 329
rect 513 322 537 326
rect 513 318 517 322
rect 559 326 563 328
rect 559 324 560 326
rect 562 324 563 326
rect 512 316 517 318
rect 512 314 513 316
rect 515 314 517 316
rect 521 317 537 318
rect 521 315 523 317
rect 525 315 537 317
rect 521 314 537 315
rect 512 312 517 314
rect 513 310 517 312
rect 513 307 529 310
rect 513 306 526 307
rect 525 305 526 306
rect 528 305 529 307
rect 525 300 529 305
rect 525 298 526 300
rect 528 298 529 300
rect 525 296 529 298
rect 533 308 537 314
rect 559 318 563 324
rect 552 314 563 318
rect 585 326 589 330
rect 622 333 642 334
rect 622 331 624 333
rect 626 331 642 333
rect 622 330 642 331
rect 600 327 601 329
rect 585 322 597 326
rect 593 317 597 322
rect 593 315 594 317
rect 596 315 597 317
rect 552 308 556 314
rect 533 307 556 308
rect 533 305 552 307
rect 554 305 556 307
rect 533 304 556 305
rect 468 291 469 293
rect 471 291 472 293
rect 468 289 472 291
rect 477 295 483 296
rect 477 293 479 295
rect 481 293 483 295
rect 533 293 537 304
rect 593 303 597 315
rect 638 326 642 330
rect 662 333 682 334
rect 662 331 664 333
rect 666 331 682 333
rect 662 330 682 331
rect 653 327 654 329
rect 638 322 650 326
rect 646 317 650 322
rect 646 315 647 317
rect 649 315 650 317
rect 580 300 597 303
rect 580 298 581 300
rect 583 299 597 300
rect 583 298 584 299
rect 477 284 483 293
rect 504 292 537 293
rect 504 290 506 292
rect 508 290 537 292
rect 504 289 537 290
rect 541 293 545 295
rect 541 291 542 293
rect 544 291 545 293
rect 541 286 545 291
rect 569 293 575 294
rect 569 291 571 293
rect 573 291 575 293
rect 541 284 542 286
rect 544 284 545 286
rect 569 284 575 291
rect 580 293 584 298
rect 646 303 650 315
rect 678 326 682 330
rect 749 334 755 340
rect 693 327 694 329
rect 678 322 690 326
rect 686 317 690 322
rect 686 315 687 317
rect 689 315 690 317
rect 633 300 650 303
rect 633 298 634 300
rect 636 299 650 300
rect 636 298 637 299
rect 580 291 581 293
rect 583 291 584 293
rect 580 289 584 291
rect 589 295 595 296
rect 589 293 591 295
rect 593 293 595 295
rect 589 284 595 293
rect 622 293 628 294
rect 622 291 624 293
rect 626 291 628 293
rect 622 284 628 291
rect 633 293 637 298
rect 686 303 690 315
rect 673 300 690 303
rect 673 298 674 300
rect 676 299 690 300
rect 676 298 677 299
rect 633 291 634 293
rect 636 291 637 293
rect 633 289 637 291
rect 642 295 648 296
rect 642 293 644 295
rect 646 293 648 295
rect 642 284 648 293
rect 662 293 668 294
rect 662 291 664 293
rect 666 291 668 293
rect 662 284 668 291
rect 673 293 677 298
rect 738 331 742 333
rect 749 332 751 334
rect 753 332 755 334
rect 749 331 755 332
rect 774 333 794 334
rect 774 331 776 333
rect 778 331 794 333
rect 738 329 739 331
rect 741 329 742 331
rect 774 330 794 331
rect 738 326 742 329
rect 718 322 742 326
rect 718 318 722 322
rect 764 326 768 328
rect 764 324 765 326
rect 767 324 768 326
rect 717 316 722 318
rect 717 314 718 316
rect 720 314 722 316
rect 726 317 742 318
rect 726 315 728 317
rect 730 315 742 317
rect 726 314 742 315
rect 717 312 722 314
rect 718 310 722 312
rect 718 307 734 310
rect 718 306 731 307
rect 730 305 731 306
rect 733 305 734 307
rect 730 300 734 305
rect 730 298 731 300
rect 733 298 734 300
rect 730 296 734 298
rect 738 308 742 314
rect 764 318 768 324
rect 757 314 768 318
rect 790 326 794 330
rect 841 333 861 334
rect 841 331 843 333
rect 845 331 861 333
rect 841 330 861 331
rect 805 327 806 329
rect 790 322 802 326
rect 798 317 802 322
rect 798 315 799 317
rect 801 315 802 317
rect 757 308 761 314
rect 738 307 761 308
rect 738 305 757 307
rect 759 305 761 307
rect 738 304 761 305
rect 673 291 674 293
rect 676 291 677 293
rect 673 289 677 291
rect 682 295 688 296
rect 682 293 684 295
rect 686 293 688 295
rect 738 293 742 304
rect 798 303 802 315
rect 857 326 861 330
rect 881 333 901 334
rect 881 331 883 333
rect 885 331 901 333
rect 881 330 901 331
rect 872 327 873 329
rect 857 322 869 326
rect 865 317 869 322
rect 865 315 866 317
rect 868 315 869 317
rect 785 300 802 303
rect 785 298 786 300
rect 788 299 802 300
rect 788 298 789 299
rect 682 284 688 293
rect 709 292 742 293
rect 709 290 711 292
rect 713 290 742 292
rect 709 289 742 290
rect 746 293 750 295
rect 746 291 747 293
rect 749 291 750 293
rect 746 286 750 291
rect 774 293 780 294
rect 774 291 776 293
rect 778 291 780 293
rect 746 284 747 286
rect 749 284 750 286
rect 774 284 780 291
rect 785 293 789 298
rect 865 303 869 315
rect 897 326 901 330
rect 968 334 974 340
rect 912 327 913 329
rect 897 322 909 326
rect 905 317 909 322
rect 905 315 906 317
rect 908 315 909 317
rect 852 300 869 303
rect 852 298 853 300
rect 855 299 869 300
rect 855 298 856 299
rect 785 291 786 293
rect 788 291 789 293
rect 785 289 789 291
rect 794 295 800 296
rect 794 293 796 295
rect 798 293 800 295
rect 794 284 800 293
rect 841 293 847 294
rect 841 291 843 293
rect 845 291 847 293
rect 841 284 847 291
rect 852 293 856 298
rect 905 303 909 315
rect 892 300 909 303
rect 892 298 893 300
rect 895 299 909 300
rect 895 298 896 299
rect 852 291 853 293
rect 855 291 856 293
rect 852 289 856 291
rect 861 295 867 296
rect 861 293 863 295
rect 865 293 867 295
rect 861 284 867 293
rect 881 293 887 294
rect 881 291 883 293
rect 885 291 887 293
rect 881 284 887 291
rect 892 293 896 298
rect 957 331 961 333
rect 968 332 970 334
rect 972 332 974 334
rect 968 331 974 332
rect 993 333 1013 334
rect 993 331 995 333
rect 997 331 1013 333
rect 957 329 958 331
rect 960 329 961 331
rect 993 330 1013 331
rect 957 326 961 329
rect 937 322 961 326
rect 937 318 941 322
rect 983 326 987 328
rect 983 324 984 326
rect 986 324 987 326
rect 936 316 941 318
rect 936 314 937 316
rect 939 314 941 316
rect 945 317 961 318
rect 945 315 947 317
rect 949 315 961 317
rect 945 314 961 315
rect 936 312 941 314
rect 937 310 941 312
rect 937 307 953 310
rect 937 306 950 307
rect 949 305 950 306
rect 952 305 953 307
rect 949 300 953 305
rect 949 298 950 300
rect 952 298 953 300
rect 949 296 953 298
rect 957 308 961 314
rect 983 318 987 324
rect 976 314 987 318
rect 1009 326 1013 330
rect 1024 327 1025 329
rect 1009 322 1021 326
rect 1017 317 1021 322
rect 1017 315 1018 317
rect 1020 315 1021 317
rect 976 308 980 314
rect 957 307 980 308
rect 957 305 976 307
rect 978 305 980 307
rect 957 304 980 305
rect 892 291 893 293
rect 895 291 896 293
rect 892 289 896 291
rect 901 295 907 296
rect 901 293 903 295
rect 905 293 907 295
rect 957 293 961 304
rect 1017 303 1021 315
rect 1004 300 1021 303
rect 1004 298 1005 300
rect 1007 299 1021 300
rect 1007 298 1008 299
rect 901 284 907 293
rect 928 292 961 293
rect 928 290 930 292
rect 932 290 961 292
rect 928 289 961 290
rect 965 293 969 295
rect 965 291 966 293
rect 968 291 969 293
rect 965 286 969 291
rect 993 293 999 294
rect 993 291 995 293
rect 997 291 999 293
rect 965 284 966 286
rect 968 284 969 286
rect 993 284 999 291
rect 1004 293 1008 298
rect 1004 291 1005 293
rect 1007 291 1008 293
rect 1004 289 1008 291
rect 1013 295 1019 296
rect 1013 293 1015 295
rect 1017 293 1019 295
rect 1013 284 1019 293
rect 211 259 217 268
rect 211 257 213 259
rect 215 257 217 259
rect 211 256 217 257
rect 222 261 226 263
rect 222 259 223 261
rect 225 259 226 261
rect 222 254 226 259
rect 231 261 237 268
rect 231 259 233 261
rect 235 259 237 261
rect 231 258 237 259
rect 241 261 247 268
rect 241 259 243 261
rect 245 259 247 261
rect 241 258 247 259
rect 252 261 256 263
rect 252 259 253 261
rect 255 259 256 261
rect 222 253 223 254
rect 209 252 223 253
rect 225 252 226 254
rect 209 249 226 252
rect 209 237 213 249
rect 252 254 256 259
rect 261 259 267 268
rect 261 257 263 259
rect 265 257 267 259
rect 261 256 267 257
rect 291 259 297 268
rect 291 257 293 259
rect 295 257 297 259
rect 291 256 297 257
rect 302 261 306 263
rect 302 259 303 261
rect 305 259 306 261
rect 252 252 253 254
rect 255 253 256 254
rect 255 252 269 253
rect 252 249 269 252
rect 209 235 210 237
rect 212 235 213 237
rect 209 230 213 235
rect 209 226 221 230
rect 205 223 206 225
rect 217 222 221 226
rect 265 237 269 249
rect 265 235 266 237
rect 268 235 269 237
rect 265 230 269 235
rect 257 226 269 230
rect 257 222 261 226
rect 272 223 273 225
rect 217 221 237 222
rect 217 219 233 221
rect 235 219 237 221
rect 217 218 237 219
rect 241 221 261 222
rect 241 219 243 221
rect 245 219 261 221
rect 241 218 261 219
rect 302 254 306 259
rect 311 261 317 268
rect 341 266 342 268
rect 344 266 345 268
rect 311 259 313 261
rect 315 259 317 261
rect 311 258 317 259
rect 341 261 345 266
rect 341 259 342 261
rect 344 259 345 261
rect 341 257 345 259
rect 349 262 382 263
rect 349 260 378 262
rect 380 260 382 262
rect 349 259 382 260
rect 427 259 433 268
rect 302 253 303 254
rect 289 252 303 253
rect 305 252 306 254
rect 289 249 306 252
rect 289 237 293 249
rect 349 248 353 259
rect 427 257 429 259
rect 431 257 433 259
rect 427 256 433 257
rect 438 261 442 263
rect 438 259 439 261
rect 441 259 442 261
rect 330 247 353 248
rect 330 245 332 247
rect 334 245 353 247
rect 330 244 353 245
rect 330 238 334 244
rect 289 235 290 237
rect 292 235 293 237
rect 289 230 293 235
rect 289 226 301 230
rect 285 223 286 225
rect 297 222 301 226
rect 323 234 334 238
rect 323 228 327 234
rect 349 238 353 244
rect 357 254 361 256
rect 357 252 358 254
rect 360 252 361 254
rect 357 247 361 252
rect 357 245 358 247
rect 360 246 361 247
rect 360 245 373 246
rect 357 242 373 245
rect 369 240 373 242
rect 369 238 374 240
rect 349 237 365 238
rect 349 235 361 237
rect 363 235 365 237
rect 349 234 365 235
rect 369 236 371 238
rect 373 236 374 238
rect 369 234 374 236
rect 323 226 324 228
rect 326 226 327 228
rect 323 224 327 226
rect 369 230 373 234
rect 349 226 373 230
rect 349 223 353 226
rect 297 221 317 222
rect 349 221 350 223
rect 352 221 353 223
rect 297 219 313 221
rect 315 219 317 221
rect 297 218 317 219
rect 336 220 342 221
rect 336 218 338 220
rect 340 218 342 220
rect 349 219 353 221
rect 438 254 442 259
rect 447 261 453 268
rect 447 259 449 261
rect 451 259 453 261
rect 447 258 453 259
rect 457 261 463 268
rect 457 259 459 261
rect 461 259 463 261
rect 457 258 463 259
rect 468 261 472 263
rect 468 259 469 261
rect 471 259 472 261
rect 438 253 439 254
rect 425 252 439 253
rect 441 252 442 254
rect 425 249 442 252
rect 425 237 429 249
rect 468 254 472 259
rect 477 259 483 268
rect 477 257 479 259
rect 481 257 483 259
rect 477 256 483 257
rect 507 259 513 268
rect 507 257 509 259
rect 511 257 513 259
rect 507 256 513 257
rect 518 261 522 263
rect 518 259 519 261
rect 521 259 522 261
rect 468 252 469 254
rect 471 253 472 254
rect 471 252 485 253
rect 468 249 485 252
rect 425 235 426 237
rect 428 235 429 237
rect 425 230 429 235
rect 425 226 437 230
rect 421 223 422 225
rect 336 212 342 218
rect 433 222 437 226
rect 481 237 485 249
rect 481 235 482 237
rect 484 235 485 237
rect 481 230 485 235
rect 473 226 485 230
rect 473 222 477 226
rect 488 223 489 225
rect 433 221 453 222
rect 433 219 449 221
rect 451 219 453 221
rect 433 218 453 219
rect 457 221 477 222
rect 457 219 459 221
rect 461 219 477 221
rect 457 218 477 219
rect 518 254 522 259
rect 527 261 533 268
rect 557 266 558 268
rect 560 266 561 268
rect 527 259 529 261
rect 531 259 533 261
rect 527 258 533 259
rect 557 261 561 266
rect 557 259 558 261
rect 560 259 561 261
rect 557 257 561 259
rect 565 262 598 263
rect 565 260 594 262
rect 596 260 598 262
rect 565 259 598 260
rect 632 259 638 268
rect 518 253 519 254
rect 505 252 519 253
rect 521 252 522 254
rect 505 249 522 252
rect 505 237 509 249
rect 565 248 569 259
rect 632 257 634 259
rect 636 257 638 259
rect 632 256 638 257
rect 643 261 647 263
rect 643 259 644 261
rect 646 259 647 261
rect 546 247 569 248
rect 546 245 548 247
rect 550 245 569 247
rect 546 244 569 245
rect 546 238 550 244
rect 505 235 506 237
rect 508 235 509 237
rect 505 230 509 235
rect 505 226 517 230
rect 501 223 502 225
rect 513 222 517 226
rect 539 234 550 238
rect 539 228 543 234
rect 565 238 569 244
rect 573 254 577 256
rect 573 252 574 254
rect 576 252 577 254
rect 573 247 577 252
rect 573 245 574 247
rect 576 246 577 247
rect 576 245 589 246
rect 573 242 589 245
rect 585 240 589 242
rect 585 238 590 240
rect 565 237 581 238
rect 565 235 577 237
rect 579 235 581 237
rect 565 234 581 235
rect 585 236 587 238
rect 589 236 590 238
rect 585 234 590 236
rect 539 226 540 228
rect 542 226 543 228
rect 539 224 543 226
rect 585 230 589 234
rect 565 226 589 230
rect 565 223 569 226
rect 513 221 533 222
rect 565 221 566 223
rect 568 221 569 223
rect 513 219 529 221
rect 531 219 533 221
rect 513 218 533 219
rect 552 220 558 221
rect 552 218 554 220
rect 556 218 558 220
rect 565 219 569 221
rect 643 254 647 259
rect 652 261 658 268
rect 652 259 654 261
rect 656 259 658 261
rect 652 258 658 259
rect 662 261 668 268
rect 662 259 664 261
rect 666 259 668 261
rect 662 258 668 259
rect 673 261 677 263
rect 673 259 674 261
rect 676 259 677 261
rect 643 253 644 254
rect 630 252 644 253
rect 646 252 647 254
rect 630 249 647 252
rect 630 237 634 249
rect 673 254 677 259
rect 682 259 688 268
rect 682 257 684 259
rect 686 257 688 259
rect 682 256 688 257
rect 712 259 718 268
rect 712 257 714 259
rect 716 257 718 259
rect 712 256 718 257
rect 723 261 727 263
rect 723 259 724 261
rect 726 259 727 261
rect 673 252 674 254
rect 676 253 677 254
rect 676 252 690 253
rect 673 249 690 252
rect 630 235 631 237
rect 633 235 634 237
rect 630 230 634 235
rect 630 226 642 230
rect 626 223 627 225
rect 552 212 558 218
rect 638 222 642 226
rect 686 237 690 249
rect 686 235 687 237
rect 689 235 690 237
rect 686 230 690 235
rect 678 226 690 230
rect 678 222 682 226
rect 693 223 694 225
rect 638 221 658 222
rect 638 219 654 221
rect 656 219 658 221
rect 638 218 658 219
rect 662 221 682 222
rect 662 219 664 221
rect 666 219 682 221
rect 662 218 682 219
rect 723 254 727 259
rect 732 261 738 268
rect 762 266 763 268
rect 765 266 766 268
rect 732 259 734 261
rect 736 259 738 261
rect 732 258 738 259
rect 762 261 766 266
rect 762 259 763 261
rect 765 259 766 261
rect 762 257 766 259
rect 770 262 803 263
rect 770 260 799 262
rect 801 260 803 262
rect 770 259 803 260
rect 851 259 857 268
rect 723 253 724 254
rect 710 252 724 253
rect 726 252 727 254
rect 710 249 727 252
rect 710 237 714 249
rect 770 248 774 259
rect 851 257 853 259
rect 855 257 857 259
rect 851 256 857 257
rect 862 261 866 263
rect 862 259 863 261
rect 865 259 866 261
rect 751 247 774 248
rect 751 245 753 247
rect 755 245 774 247
rect 751 244 774 245
rect 751 238 755 244
rect 710 235 711 237
rect 713 235 714 237
rect 710 230 714 235
rect 710 226 722 230
rect 706 223 707 225
rect 718 222 722 226
rect 744 234 755 238
rect 744 228 748 234
rect 770 238 774 244
rect 778 254 782 256
rect 778 252 779 254
rect 781 252 782 254
rect 778 247 782 252
rect 778 245 779 247
rect 781 246 782 247
rect 781 245 794 246
rect 778 242 794 245
rect 790 240 794 242
rect 790 238 795 240
rect 770 237 786 238
rect 770 235 782 237
rect 784 235 786 237
rect 770 234 786 235
rect 790 236 792 238
rect 794 236 795 238
rect 790 234 795 236
rect 744 226 745 228
rect 747 226 748 228
rect 744 224 748 226
rect 790 230 794 234
rect 770 226 794 230
rect 770 223 774 226
rect 718 221 738 222
rect 770 221 771 223
rect 773 221 774 223
rect 718 219 734 221
rect 736 219 738 221
rect 718 218 738 219
rect 757 220 763 221
rect 757 218 759 220
rect 761 218 763 220
rect 770 219 774 221
rect 862 254 866 259
rect 871 261 877 268
rect 871 259 873 261
rect 875 259 877 261
rect 871 258 877 259
rect 881 261 887 268
rect 881 259 883 261
rect 885 259 887 261
rect 881 258 887 259
rect 892 261 896 263
rect 892 259 893 261
rect 895 259 896 261
rect 862 253 863 254
rect 849 252 863 253
rect 865 252 866 254
rect 849 249 866 252
rect 849 237 853 249
rect 892 254 896 259
rect 901 259 907 268
rect 901 257 903 259
rect 905 257 907 259
rect 901 256 907 257
rect 931 259 937 268
rect 931 257 933 259
rect 935 257 937 259
rect 931 256 937 257
rect 942 261 946 263
rect 942 259 943 261
rect 945 259 946 261
rect 892 252 893 254
rect 895 253 896 254
rect 895 252 909 253
rect 892 249 909 252
rect 849 235 850 237
rect 852 235 853 237
rect 849 230 853 235
rect 849 226 861 230
rect 845 223 846 225
rect 757 212 763 218
rect 857 222 861 226
rect 905 237 909 249
rect 905 235 906 237
rect 908 235 909 237
rect 905 230 909 235
rect 897 226 909 230
rect 897 222 901 226
rect 912 223 913 225
rect 857 221 877 222
rect 857 219 873 221
rect 875 219 877 221
rect 857 218 877 219
rect 881 221 901 222
rect 881 219 883 221
rect 885 219 901 221
rect 881 218 901 219
rect 942 254 946 259
rect 951 261 957 268
rect 981 266 982 268
rect 984 266 985 268
rect 951 259 953 261
rect 955 259 957 261
rect 951 258 957 259
rect 981 261 985 266
rect 981 259 982 261
rect 984 259 985 261
rect 981 257 985 259
rect 989 262 1022 263
rect 989 260 1018 262
rect 1020 260 1022 262
rect 989 259 1022 260
rect 1055 259 1061 268
rect 942 253 943 254
rect 929 252 943 253
rect 945 252 946 254
rect 929 249 946 252
rect 929 237 933 249
rect 989 248 993 259
rect 1055 257 1057 259
rect 1059 257 1061 259
rect 1055 256 1061 257
rect 1066 261 1070 263
rect 1066 259 1067 261
rect 1069 259 1070 261
rect 970 247 993 248
rect 970 245 972 247
rect 974 245 993 247
rect 970 244 993 245
rect 970 238 974 244
rect 929 235 930 237
rect 932 235 933 237
rect 929 230 933 235
rect 929 226 941 230
rect 925 223 926 225
rect 937 222 941 226
rect 963 234 974 238
rect 963 228 967 234
rect 989 238 993 244
rect 997 254 1001 256
rect 997 252 998 254
rect 1000 252 1001 254
rect 997 247 1001 252
rect 997 245 998 247
rect 1000 246 1001 247
rect 1000 245 1013 246
rect 997 242 1013 245
rect 1009 240 1013 242
rect 1009 238 1014 240
rect 989 237 1005 238
rect 989 235 1001 237
rect 1003 235 1005 237
rect 989 234 1005 235
rect 1009 236 1011 238
rect 1013 236 1014 238
rect 1009 234 1014 236
rect 963 226 964 228
rect 966 226 967 228
rect 963 224 967 226
rect 1009 230 1013 234
rect 989 226 1013 230
rect 989 223 993 226
rect 937 221 957 222
rect 989 221 990 223
rect 992 221 993 223
rect 937 219 953 221
rect 955 219 957 221
rect 937 218 957 219
rect 976 220 982 221
rect 976 218 978 220
rect 980 218 982 220
rect 989 219 993 221
rect 1066 254 1070 259
rect 1075 261 1081 268
rect 1105 266 1106 268
rect 1108 266 1109 268
rect 1075 259 1077 261
rect 1079 259 1081 261
rect 1075 258 1081 259
rect 1105 261 1109 266
rect 1105 259 1106 261
rect 1108 259 1109 261
rect 1105 257 1109 259
rect 1113 262 1146 263
rect 1113 260 1142 262
rect 1144 260 1146 262
rect 1113 259 1146 260
rect 1066 253 1067 254
rect 1053 252 1067 253
rect 1069 252 1070 254
rect 1053 249 1070 252
rect 1053 237 1057 249
rect 1113 248 1117 259
rect 1094 247 1117 248
rect 1094 245 1096 247
rect 1098 245 1117 247
rect 1094 244 1117 245
rect 1094 238 1098 244
rect 1053 235 1054 237
rect 1056 235 1057 237
rect 1053 230 1057 235
rect 1053 226 1065 230
rect 1049 223 1050 225
rect 976 212 982 218
rect 1061 222 1065 226
rect 1087 234 1098 238
rect 1087 228 1091 234
rect 1113 238 1117 244
rect 1121 254 1125 256
rect 1121 252 1122 254
rect 1124 252 1125 254
rect 1121 247 1125 252
rect 1121 245 1122 247
rect 1124 246 1125 247
rect 1124 245 1137 246
rect 1121 242 1137 245
rect 1133 240 1137 242
rect 1133 238 1138 240
rect 1113 237 1129 238
rect 1113 235 1125 237
rect 1127 235 1129 237
rect 1113 234 1129 235
rect 1133 236 1135 238
rect 1137 236 1138 238
rect 1133 234 1138 236
rect 1087 226 1088 228
rect 1090 226 1091 228
rect 1087 224 1091 226
rect 1133 230 1137 234
rect 1113 226 1137 230
rect 1113 223 1117 226
rect 1061 221 1081 222
rect 1113 221 1114 223
rect 1116 221 1117 223
rect 1061 219 1077 221
rect 1079 219 1081 221
rect 1061 218 1081 219
rect 1100 220 1106 221
rect 1100 218 1102 220
rect 1104 218 1106 220
rect 1113 219 1117 221
rect 1100 212 1106 218
rect 162 195 168 196
rect 162 193 164 195
rect 166 193 168 195
rect 162 192 168 193
rect 181 195 187 196
rect 181 193 183 195
rect 185 193 187 195
rect 181 192 187 193
rect 246 190 252 196
rect 207 189 227 190
rect 207 187 223 189
rect 225 187 227 189
rect 246 188 248 190
rect 250 188 252 190
rect 246 187 252 188
rect 259 187 263 189
rect 207 186 227 187
rect 159 182 177 183
rect 159 180 173 182
rect 175 180 177 182
rect 159 179 177 180
rect 159 173 163 179
rect 195 183 196 185
rect 207 182 211 186
rect 259 185 260 187
rect 262 185 263 187
rect 159 171 160 173
rect 162 171 163 173
rect 155 150 156 161
rect 159 158 163 171
rect 178 166 184 167
rect 159 154 174 158
rect 170 150 174 154
rect 199 178 211 182
rect 199 173 203 178
rect 199 171 200 173
rect 202 171 203 173
rect 199 159 203 171
rect 233 182 237 184
rect 233 180 234 182
rect 236 180 237 182
rect 233 174 237 180
rect 259 182 263 185
rect 259 178 283 182
rect 233 170 244 174
rect 240 164 244 170
rect 279 174 283 178
rect 259 173 275 174
rect 259 171 271 173
rect 273 171 275 173
rect 259 170 275 171
rect 279 172 284 174
rect 279 170 281 172
rect 283 170 284 172
rect 259 164 263 170
rect 279 168 284 170
rect 279 166 283 168
rect 240 163 263 164
rect 240 161 242 163
rect 244 161 263 163
rect 240 160 263 161
rect 199 156 216 159
rect 199 155 213 156
rect 212 154 213 155
rect 215 154 216 156
rect 201 151 207 152
rect 170 149 187 150
rect 170 147 183 149
rect 185 147 187 149
rect 170 146 187 147
rect 201 149 203 151
rect 205 149 207 151
rect 162 142 168 143
rect 162 140 164 142
rect 166 140 168 142
rect 201 140 207 149
rect 212 149 216 154
rect 212 147 213 149
rect 215 147 216 149
rect 212 145 216 147
rect 221 149 227 150
rect 221 147 223 149
rect 225 147 227 149
rect 221 140 227 147
rect 251 149 255 151
rect 251 147 252 149
rect 254 147 255 149
rect 251 142 255 147
rect 259 149 263 160
rect 267 163 283 166
rect 267 161 268 163
rect 270 162 283 163
rect 270 161 271 162
rect 267 156 271 161
rect 267 154 268 156
rect 270 154 271 156
rect 267 152 271 154
rect 351 190 357 196
rect 412 195 418 196
rect 412 193 414 195
rect 416 193 418 195
rect 412 192 418 193
rect 431 195 437 196
rect 431 193 433 195
rect 435 193 437 195
rect 431 192 437 193
rect 312 189 332 190
rect 312 187 328 189
rect 330 187 332 189
rect 351 188 353 190
rect 355 188 357 190
rect 351 187 357 188
rect 364 187 368 189
rect 312 186 332 187
rect 300 183 301 185
rect 312 182 316 186
rect 364 185 365 187
rect 367 185 368 187
rect 304 178 316 182
rect 304 173 308 178
rect 304 171 305 173
rect 307 171 308 173
rect 304 159 308 171
rect 338 182 342 184
rect 338 180 339 182
rect 341 180 342 182
rect 338 174 342 180
rect 364 182 368 185
rect 364 178 388 182
rect 338 170 349 174
rect 345 164 349 170
rect 384 174 388 178
rect 364 173 380 174
rect 364 171 376 173
rect 378 171 380 173
rect 364 170 380 171
rect 384 172 389 174
rect 384 170 386 172
rect 388 170 389 172
rect 364 164 368 170
rect 384 168 389 170
rect 384 166 388 168
rect 345 163 368 164
rect 345 161 347 163
rect 349 161 368 163
rect 345 160 368 161
rect 304 156 321 159
rect 304 155 318 156
rect 317 154 318 155
rect 320 154 321 156
rect 306 151 312 152
rect 306 149 308 151
rect 310 149 312 151
rect 259 148 292 149
rect 259 146 288 148
rect 290 146 292 148
rect 259 145 292 146
rect 251 140 252 142
rect 254 140 255 142
rect 306 140 312 149
rect 317 149 321 154
rect 317 147 318 149
rect 320 147 321 149
rect 317 145 321 147
rect 326 149 332 150
rect 326 147 328 149
rect 330 147 332 149
rect 326 140 332 147
rect 356 149 360 151
rect 356 147 357 149
rect 359 147 360 149
rect 356 142 360 147
rect 364 149 368 160
rect 372 163 388 166
rect 372 161 373 163
rect 375 162 388 163
rect 375 161 376 162
rect 372 156 376 161
rect 496 190 502 196
rect 457 189 477 190
rect 457 187 473 189
rect 475 187 477 189
rect 496 188 498 190
rect 500 188 502 190
rect 496 187 502 188
rect 509 187 513 189
rect 457 186 477 187
rect 372 154 373 156
rect 375 154 376 156
rect 372 152 376 154
rect 409 182 427 183
rect 409 180 423 182
rect 425 180 427 182
rect 409 179 427 180
rect 409 173 413 179
rect 445 183 446 185
rect 457 182 461 186
rect 509 185 510 187
rect 512 185 513 187
rect 409 171 410 173
rect 412 171 413 173
rect 405 150 406 161
rect 409 158 413 171
rect 428 166 434 167
rect 409 154 424 158
rect 420 150 424 154
rect 449 178 461 182
rect 449 173 453 178
rect 449 171 450 173
rect 452 171 453 173
rect 449 159 453 171
rect 483 182 487 184
rect 483 180 484 182
rect 486 180 487 182
rect 483 174 487 180
rect 509 182 513 185
rect 509 178 533 182
rect 483 170 494 174
rect 490 164 494 170
rect 529 174 533 178
rect 509 173 525 174
rect 509 171 521 173
rect 523 171 525 173
rect 509 170 525 171
rect 529 172 534 174
rect 529 170 531 172
rect 533 170 534 172
rect 509 164 513 170
rect 529 168 534 170
rect 529 166 533 168
rect 490 163 513 164
rect 490 161 492 163
rect 494 161 513 163
rect 490 160 513 161
rect 449 156 466 159
rect 449 155 463 156
rect 462 154 463 155
rect 465 154 466 156
rect 451 151 457 152
rect 364 148 397 149
rect 364 146 393 148
rect 395 146 397 148
rect 364 145 397 146
rect 420 149 437 150
rect 420 147 433 149
rect 435 147 437 149
rect 420 146 437 147
rect 451 149 453 151
rect 455 149 457 151
rect 356 140 357 142
rect 359 140 360 142
rect 412 142 418 143
rect 412 140 414 142
rect 416 140 418 142
rect 451 140 457 149
rect 462 149 466 154
rect 462 147 463 149
rect 465 147 466 149
rect 462 145 466 147
rect 471 149 477 150
rect 471 147 473 149
rect 475 147 477 149
rect 471 140 477 147
rect 501 149 505 151
rect 501 147 502 149
rect 504 147 505 149
rect 501 142 505 147
rect 509 149 513 160
rect 517 163 533 166
rect 517 161 518 163
rect 520 162 533 163
rect 520 161 521 162
rect 517 156 521 161
rect 517 154 518 156
rect 520 154 521 156
rect 517 152 521 154
rect 601 190 607 196
rect 662 195 668 196
rect 662 193 664 195
rect 666 193 668 195
rect 662 192 668 193
rect 681 195 687 196
rect 681 193 683 195
rect 685 193 687 195
rect 681 192 687 193
rect 562 189 582 190
rect 562 187 578 189
rect 580 187 582 189
rect 601 188 603 190
rect 605 188 607 190
rect 601 187 607 188
rect 614 187 618 189
rect 562 186 582 187
rect 550 183 551 185
rect 562 182 566 186
rect 614 185 615 187
rect 617 185 618 187
rect 554 178 566 182
rect 554 173 558 178
rect 554 171 555 173
rect 557 171 558 173
rect 554 159 558 171
rect 588 182 592 184
rect 588 180 589 182
rect 591 180 592 182
rect 588 174 592 180
rect 614 182 618 185
rect 614 178 638 182
rect 588 170 599 174
rect 595 164 599 170
rect 634 174 638 178
rect 614 173 630 174
rect 614 171 626 173
rect 628 171 630 173
rect 614 170 630 171
rect 634 172 639 174
rect 634 170 636 172
rect 638 170 639 172
rect 614 164 618 170
rect 634 168 639 170
rect 634 166 638 168
rect 595 163 618 164
rect 595 161 597 163
rect 599 161 618 163
rect 595 160 618 161
rect 554 156 571 159
rect 554 155 568 156
rect 567 154 568 155
rect 570 154 571 156
rect 556 151 562 152
rect 556 149 558 151
rect 560 149 562 151
rect 509 148 542 149
rect 509 146 538 148
rect 540 146 542 148
rect 509 145 542 146
rect 501 140 502 142
rect 504 140 505 142
rect 556 140 562 149
rect 567 149 571 154
rect 567 147 568 149
rect 570 147 571 149
rect 567 145 571 147
rect 576 149 582 150
rect 576 147 578 149
rect 580 147 582 149
rect 576 140 582 147
rect 606 149 610 151
rect 606 147 607 149
rect 609 147 610 149
rect 606 142 610 147
rect 614 149 618 160
rect 622 163 638 166
rect 622 161 623 163
rect 625 162 638 163
rect 625 161 626 162
rect 622 156 626 161
rect 746 190 752 196
rect 707 189 727 190
rect 707 187 723 189
rect 725 187 727 189
rect 746 188 748 190
rect 750 188 752 190
rect 746 187 752 188
rect 759 187 763 189
rect 707 186 727 187
rect 622 154 623 156
rect 625 154 626 156
rect 622 152 626 154
rect 659 182 677 183
rect 659 180 673 182
rect 675 180 677 182
rect 659 179 677 180
rect 659 173 663 179
rect 695 183 696 185
rect 707 182 711 186
rect 759 185 760 187
rect 762 185 763 187
rect 659 171 660 173
rect 662 171 663 173
rect 655 150 656 161
rect 659 158 663 171
rect 678 166 684 167
rect 659 154 674 158
rect 670 150 674 154
rect 699 178 711 182
rect 699 173 703 178
rect 699 171 700 173
rect 702 171 703 173
rect 699 159 703 171
rect 733 182 737 184
rect 733 180 734 182
rect 736 180 737 182
rect 733 174 737 180
rect 759 182 763 185
rect 759 178 783 182
rect 733 170 744 174
rect 740 164 744 170
rect 779 174 783 178
rect 759 173 775 174
rect 759 171 771 173
rect 773 171 775 173
rect 759 170 775 171
rect 779 172 784 174
rect 779 170 781 172
rect 783 170 784 172
rect 759 164 763 170
rect 779 168 784 170
rect 779 166 783 168
rect 740 163 763 164
rect 740 161 742 163
rect 744 161 763 163
rect 740 160 763 161
rect 699 156 716 159
rect 699 155 713 156
rect 712 154 713 155
rect 715 154 716 156
rect 701 151 707 152
rect 614 148 647 149
rect 614 146 643 148
rect 645 146 647 148
rect 614 145 647 146
rect 670 149 687 150
rect 670 147 683 149
rect 685 147 687 149
rect 670 146 687 147
rect 701 149 703 151
rect 705 149 707 151
rect 606 140 607 142
rect 609 140 610 142
rect 662 142 668 143
rect 662 140 664 142
rect 666 140 668 142
rect 701 140 707 149
rect 712 149 716 154
rect 712 147 713 149
rect 715 147 716 149
rect 712 145 716 147
rect 721 149 727 150
rect 721 147 723 149
rect 725 147 727 149
rect 721 140 727 147
rect 751 149 755 151
rect 751 147 752 149
rect 754 147 755 149
rect 751 142 755 147
rect 759 149 763 160
rect 767 163 783 166
rect 767 161 768 163
rect 770 162 783 163
rect 770 161 771 162
rect 767 156 771 161
rect 767 154 768 156
rect 770 154 771 156
rect 767 152 771 154
rect 851 190 857 196
rect 912 195 918 196
rect 912 193 914 195
rect 916 193 918 195
rect 912 192 918 193
rect 931 195 937 196
rect 931 193 933 195
rect 935 193 937 195
rect 931 192 937 193
rect 812 189 832 190
rect 812 187 828 189
rect 830 187 832 189
rect 851 188 853 190
rect 855 188 857 190
rect 851 187 857 188
rect 864 187 868 189
rect 812 186 832 187
rect 800 183 801 185
rect 812 182 816 186
rect 864 185 865 187
rect 867 185 868 187
rect 804 178 816 182
rect 804 173 808 178
rect 804 171 805 173
rect 807 171 808 173
rect 804 159 808 171
rect 838 182 842 184
rect 838 180 839 182
rect 841 180 842 182
rect 838 174 842 180
rect 864 182 868 185
rect 864 178 888 182
rect 838 170 849 174
rect 845 164 849 170
rect 884 174 888 178
rect 864 173 880 174
rect 864 171 876 173
rect 878 171 880 173
rect 864 170 880 171
rect 884 172 889 174
rect 884 170 886 172
rect 888 170 889 172
rect 864 164 868 170
rect 884 168 889 170
rect 884 166 888 168
rect 845 163 868 164
rect 845 161 847 163
rect 849 161 868 163
rect 845 160 868 161
rect 804 156 821 159
rect 804 155 818 156
rect 817 154 818 155
rect 820 154 821 156
rect 806 151 812 152
rect 806 149 808 151
rect 810 149 812 151
rect 759 148 792 149
rect 759 146 788 148
rect 790 146 792 148
rect 759 145 792 146
rect 751 140 752 142
rect 754 140 755 142
rect 806 140 812 149
rect 817 149 821 154
rect 817 147 818 149
rect 820 147 821 149
rect 817 145 821 147
rect 826 149 832 150
rect 826 147 828 149
rect 830 147 832 149
rect 826 140 832 147
rect 856 149 860 151
rect 856 147 857 149
rect 859 147 860 149
rect 856 142 860 147
rect 864 149 868 160
rect 872 163 888 166
rect 872 161 873 163
rect 875 162 888 163
rect 875 161 876 162
rect 872 156 876 161
rect 996 190 1002 196
rect 957 189 977 190
rect 957 187 973 189
rect 975 187 977 189
rect 996 188 998 190
rect 1000 188 1002 190
rect 996 187 1002 188
rect 1009 187 1013 189
rect 957 186 977 187
rect 872 154 873 156
rect 875 154 876 156
rect 872 152 876 154
rect 909 182 927 183
rect 909 180 923 182
rect 925 180 927 182
rect 909 179 927 180
rect 909 173 913 179
rect 945 183 946 185
rect 957 182 961 186
rect 1009 185 1010 187
rect 1012 185 1013 187
rect 909 171 910 173
rect 912 171 913 173
rect 905 150 906 161
rect 909 158 913 171
rect 928 166 934 167
rect 909 154 924 158
rect 920 150 924 154
rect 949 178 961 182
rect 949 173 953 178
rect 949 171 950 173
rect 952 171 953 173
rect 949 159 953 171
rect 983 182 987 184
rect 983 180 984 182
rect 986 180 987 182
rect 983 174 987 180
rect 1009 182 1013 185
rect 1009 178 1033 182
rect 983 170 994 174
rect 990 164 994 170
rect 1029 174 1033 178
rect 1009 173 1025 174
rect 1009 171 1021 173
rect 1023 171 1025 173
rect 1009 170 1025 171
rect 1029 172 1034 174
rect 1029 170 1031 172
rect 1033 170 1034 172
rect 1009 164 1013 170
rect 1029 168 1034 170
rect 1029 166 1033 168
rect 990 163 1013 164
rect 990 161 992 163
rect 994 161 1013 163
rect 990 160 1013 161
rect 949 156 966 159
rect 949 155 963 156
rect 962 154 963 155
rect 965 154 966 156
rect 951 151 957 152
rect 864 148 897 149
rect 864 146 893 148
rect 895 146 897 148
rect 864 145 897 146
rect 920 149 937 150
rect 920 147 933 149
rect 935 147 937 149
rect 920 146 937 147
rect 951 149 953 151
rect 955 149 957 151
rect 856 140 857 142
rect 859 140 860 142
rect 912 142 918 143
rect 912 140 914 142
rect 916 140 918 142
rect 951 140 957 149
rect 962 149 966 154
rect 962 147 963 149
rect 965 147 966 149
rect 962 145 966 147
rect 971 149 977 150
rect 971 147 973 149
rect 975 147 977 149
rect 971 140 977 147
rect 1001 149 1005 151
rect 1001 147 1002 149
rect 1004 147 1005 149
rect 1001 142 1005 147
rect 1009 149 1013 160
rect 1017 163 1033 166
rect 1017 161 1018 163
rect 1020 162 1033 163
rect 1020 161 1021 162
rect 1017 156 1021 161
rect 1017 154 1018 156
rect 1020 154 1021 156
rect 1017 152 1021 154
rect 1101 190 1107 196
rect 1062 189 1082 190
rect 1062 187 1078 189
rect 1080 187 1082 189
rect 1101 188 1103 190
rect 1105 188 1107 190
rect 1101 187 1107 188
rect 1114 187 1118 189
rect 1062 186 1082 187
rect 1050 183 1051 185
rect 1062 182 1066 186
rect 1114 185 1115 187
rect 1117 185 1118 187
rect 1054 178 1066 182
rect 1054 173 1058 178
rect 1054 171 1055 173
rect 1057 171 1058 173
rect 1054 159 1058 171
rect 1088 182 1092 184
rect 1088 180 1089 182
rect 1091 180 1092 182
rect 1088 174 1092 180
rect 1114 182 1118 185
rect 1114 178 1138 182
rect 1088 170 1099 174
rect 1095 164 1099 170
rect 1134 174 1138 178
rect 1114 173 1130 174
rect 1114 171 1126 173
rect 1128 171 1130 173
rect 1114 170 1130 171
rect 1134 172 1139 174
rect 1134 170 1136 172
rect 1138 170 1139 172
rect 1114 164 1118 170
rect 1134 168 1139 170
rect 1134 166 1138 168
rect 1095 163 1118 164
rect 1095 161 1097 163
rect 1099 161 1118 163
rect 1095 160 1118 161
rect 1054 156 1071 159
rect 1054 155 1068 156
rect 1067 154 1068 155
rect 1070 154 1071 156
rect 1056 151 1062 152
rect 1056 149 1058 151
rect 1060 149 1062 151
rect 1009 148 1042 149
rect 1009 146 1038 148
rect 1040 146 1042 148
rect 1009 145 1042 146
rect 1001 140 1002 142
rect 1004 140 1005 142
rect 1056 140 1062 149
rect 1067 149 1071 154
rect 1067 147 1068 149
rect 1070 147 1071 149
rect 1067 145 1071 147
rect 1076 149 1082 150
rect 1076 147 1078 149
rect 1080 147 1082 149
rect 1076 140 1082 147
rect 1106 149 1110 151
rect 1106 147 1107 149
rect 1109 147 1110 149
rect 1106 142 1110 147
rect 1114 149 1118 160
rect 1122 163 1138 166
rect 1122 161 1123 163
rect 1125 162 1138 163
rect 1125 161 1126 162
rect 1122 156 1126 161
rect 1122 154 1123 156
rect 1125 154 1126 156
rect 1122 152 1126 154
rect 1114 148 1147 149
rect 1114 146 1143 148
rect 1145 146 1147 148
rect 1114 145 1147 146
rect 1106 140 1107 142
rect 1109 140 1110 142
rect 161 122 163 124
rect 165 122 167 124
rect 161 121 167 122
rect 169 117 186 118
rect 169 115 182 117
rect 184 115 186 117
rect 169 114 186 115
rect 200 115 206 124
rect 154 103 155 114
rect 169 110 173 114
rect 200 113 202 115
rect 204 113 206 115
rect 200 112 206 113
rect 211 117 215 119
rect 211 115 212 117
rect 214 115 215 117
rect 158 106 173 110
rect 158 93 162 106
rect 211 110 215 115
rect 220 117 226 124
rect 250 122 251 124
rect 253 122 254 124
rect 220 115 222 117
rect 224 115 226 117
rect 220 114 226 115
rect 250 117 254 122
rect 250 115 251 117
rect 253 115 254 117
rect 250 113 254 115
rect 258 118 291 119
rect 258 116 287 118
rect 289 116 291 118
rect 258 115 291 116
rect 305 115 311 124
rect 211 109 212 110
rect 198 108 212 109
rect 214 108 215 110
rect 198 105 215 108
rect 177 97 183 98
rect 158 91 159 93
rect 161 91 162 93
rect 158 85 162 91
rect 158 84 176 85
rect 158 82 172 84
rect 174 82 176 84
rect 158 81 176 82
rect 198 93 202 105
rect 258 104 262 115
rect 305 113 307 115
rect 309 113 311 115
rect 305 112 311 113
rect 316 117 320 119
rect 316 115 317 117
rect 319 115 320 117
rect 239 103 262 104
rect 239 101 241 103
rect 243 101 262 103
rect 239 100 262 101
rect 239 94 243 100
rect 198 91 199 93
rect 201 91 202 93
rect 198 86 202 91
rect 198 82 210 86
rect 194 79 195 81
rect 206 78 210 82
rect 232 90 243 94
rect 232 84 236 90
rect 258 94 262 100
rect 266 110 270 112
rect 266 108 267 110
rect 269 108 270 110
rect 266 103 270 108
rect 266 101 267 103
rect 269 102 270 103
rect 269 101 282 102
rect 266 98 282 101
rect 278 96 282 98
rect 278 94 283 96
rect 258 93 274 94
rect 258 91 270 93
rect 272 91 274 93
rect 258 90 274 91
rect 278 92 280 94
rect 282 92 283 94
rect 278 90 283 92
rect 232 82 233 84
rect 235 82 236 84
rect 232 80 236 82
rect 278 86 282 90
rect 258 82 282 86
rect 258 79 262 82
rect 206 77 226 78
rect 258 77 259 79
rect 261 77 262 79
rect 206 75 222 77
rect 224 75 226 77
rect 206 74 226 75
rect 245 76 251 77
rect 245 74 247 76
rect 249 74 251 76
rect 258 75 262 77
rect 316 110 320 115
rect 325 117 331 124
rect 355 122 356 124
rect 358 122 359 124
rect 325 115 327 117
rect 329 115 331 117
rect 325 114 331 115
rect 355 117 359 122
rect 411 122 413 124
rect 415 122 417 124
rect 411 121 417 122
rect 355 115 356 117
rect 358 115 359 117
rect 355 113 359 115
rect 363 118 396 119
rect 363 116 392 118
rect 394 116 396 118
rect 363 115 396 116
rect 316 109 317 110
rect 303 108 317 109
rect 319 108 320 110
rect 303 105 320 108
rect 303 93 307 105
rect 363 104 367 115
rect 419 117 436 118
rect 419 115 432 117
rect 434 115 436 117
rect 419 114 436 115
rect 450 115 456 124
rect 344 103 367 104
rect 344 101 346 103
rect 348 101 367 103
rect 344 100 367 101
rect 344 94 348 100
rect 303 91 304 93
rect 306 91 307 93
rect 303 86 307 91
rect 303 82 315 86
rect 299 79 300 81
rect 161 71 167 72
rect 161 69 163 71
rect 165 69 167 71
rect 161 68 167 69
rect 180 71 186 72
rect 180 69 182 71
rect 184 69 186 71
rect 180 68 186 69
rect 245 68 251 74
rect 311 78 315 82
rect 337 90 348 94
rect 337 84 341 90
rect 363 94 367 100
rect 371 110 375 112
rect 371 108 372 110
rect 374 108 375 110
rect 371 103 375 108
rect 371 101 372 103
rect 374 102 375 103
rect 374 101 387 102
rect 371 98 387 101
rect 383 96 387 98
rect 383 94 388 96
rect 363 93 379 94
rect 363 91 375 93
rect 377 91 379 93
rect 363 90 379 91
rect 383 92 385 94
rect 387 92 388 94
rect 383 90 388 92
rect 337 82 338 84
rect 340 82 341 84
rect 337 80 341 82
rect 383 86 387 90
rect 363 82 387 86
rect 363 79 367 82
rect 311 77 331 78
rect 363 77 364 79
rect 366 77 367 79
rect 404 103 405 114
rect 419 110 423 114
rect 450 113 452 115
rect 454 113 456 115
rect 450 112 456 113
rect 461 117 465 119
rect 461 115 462 117
rect 464 115 465 117
rect 408 106 423 110
rect 408 93 412 106
rect 461 110 465 115
rect 470 117 476 124
rect 500 122 501 124
rect 503 122 504 124
rect 470 115 472 117
rect 474 115 476 117
rect 470 114 476 115
rect 500 117 504 122
rect 500 115 501 117
rect 503 115 504 117
rect 500 113 504 115
rect 508 118 541 119
rect 508 116 537 118
rect 539 116 541 118
rect 508 115 541 116
rect 555 115 561 124
rect 461 109 462 110
rect 448 108 462 109
rect 464 108 465 110
rect 448 105 465 108
rect 427 97 433 98
rect 408 91 409 93
rect 411 91 412 93
rect 408 85 412 91
rect 408 84 426 85
rect 408 82 422 84
rect 424 82 426 84
rect 408 81 426 82
rect 311 75 327 77
rect 329 75 331 77
rect 311 74 331 75
rect 350 76 356 77
rect 350 74 352 76
rect 354 74 356 76
rect 363 75 367 77
rect 448 93 452 105
rect 508 104 512 115
rect 555 113 557 115
rect 559 113 561 115
rect 555 112 561 113
rect 566 117 570 119
rect 566 115 567 117
rect 569 115 570 117
rect 489 103 512 104
rect 489 101 491 103
rect 493 101 512 103
rect 489 100 512 101
rect 489 94 493 100
rect 448 91 449 93
rect 451 91 452 93
rect 448 86 452 91
rect 448 82 460 86
rect 444 79 445 81
rect 350 68 356 74
rect 456 78 460 82
rect 482 90 493 94
rect 482 84 486 90
rect 508 94 512 100
rect 516 110 520 112
rect 516 108 517 110
rect 519 108 520 110
rect 516 103 520 108
rect 516 101 517 103
rect 519 102 520 103
rect 519 101 532 102
rect 516 98 532 101
rect 528 96 532 98
rect 528 94 533 96
rect 508 93 524 94
rect 508 91 520 93
rect 522 91 524 93
rect 508 90 524 91
rect 528 92 530 94
rect 532 92 533 94
rect 528 90 533 92
rect 482 82 483 84
rect 485 82 486 84
rect 482 80 486 82
rect 528 86 532 90
rect 508 82 532 86
rect 508 79 512 82
rect 456 77 476 78
rect 508 77 509 79
rect 511 77 512 79
rect 456 75 472 77
rect 474 75 476 77
rect 456 74 476 75
rect 495 76 501 77
rect 495 74 497 76
rect 499 74 501 76
rect 508 75 512 77
rect 566 110 570 115
rect 575 117 581 124
rect 605 122 606 124
rect 608 122 609 124
rect 575 115 577 117
rect 579 115 581 117
rect 575 114 581 115
rect 605 117 609 122
rect 661 122 663 124
rect 665 122 667 124
rect 661 121 667 122
rect 605 115 606 117
rect 608 115 609 117
rect 605 113 609 115
rect 613 118 646 119
rect 613 116 642 118
rect 644 116 646 118
rect 613 115 646 116
rect 566 109 567 110
rect 553 108 567 109
rect 569 108 570 110
rect 553 105 570 108
rect 553 93 557 105
rect 613 104 617 115
rect 669 117 686 118
rect 669 115 682 117
rect 684 115 686 117
rect 669 114 686 115
rect 700 115 706 124
rect 594 103 617 104
rect 594 101 596 103
rect 598 101 617 103
rect 594 100 617 101
rect 594 94 598 100
rect 553 91 554 93
rect 556 91 557 93
rect 553 86 557 91
rect 553 82 565 86
rect 549 79 550 81
rect 411 71 417 72
rect 411 69 413 71
rect 415 69 417 71
rect 411 68 417 69
rect 430 71 436 72
rect 430 69 432 71
rect 434 69 436 71
rect 430 68 436 69
rect 495 68 501 74
rect 561 78 565 82
rect 587 90 598 94
rect 587 84 591 90
rect 613 94 617 100
rect 621 110 625 112
rect 621 108 622 110
rect 624 108 625 110
rect 621 103 625 108
rect 621 101 622 103
rect 624 102 625 103
rect 624 101 637 102
rect 621 98 637 101
rect 633 96 637 98
rect 633 94 638 96
rect 613 93 629 94
rect 613 91 625 93
rect 627 91 629 93
rect 613 90 629 91
rect 633 92 635 94
rect 637 92 638 94
rect 633 90 638 92
rect 587 82 588 84
rect 590 82 591 84
rect 587 80 591 82
rect 633 86 637 90
rect 613 82 637 86
rect 613 79 617 82
rect 561 77 581 78
rect 613 77 614 79
rect 616 77 617 79
rect 654 103 655 114
rect 669 110 673 114
rect 700 113 702 115
rect 704 113 706 115
rect 700 112 706 113
rect 711 117 715 119
rect 711 115 712 117
rect 714 115 715 117
rect 658 106 673 110
rect 658 93 662 106
rect 711 110 715 115
rect 720 117 726 124
rect 750 122 751 124
rect 753 122 754 124
rect 720 115 722 117
rect 724 115 726 117
rect 720 114 726 115
rect 750 117 754 122
rect 750 115 751 117
rect 753 115 754 117
rect 750 113 754 115
rect 758 118 791 119
rect 758 116 787 118
rect 789 116 791 118
rect 758 115 791 116
rect 805 115 811 124
rect 711 109 712 110
rect 698 108 712 109
rect 714 108 715 110
rect 698 105 715 108
rect 677 97 683 98
rect 658 91 659 93
rect 661 91 662 93
rect 658 85 662 91
rect 658 84 676 85
rect 658 82 672 84
rect 674 82 676 84
rect 658 81 676 82
rect 561 75 577 77
rect 579 75 581 77
rect 561 74 581 75
rect 600 76 606 77
rect 600 74 602 76
rect 604 74 606 76
rect 613 75 617 77
rect 698 93 702 105
rect 758 104 762 115
rect 805 113 807 115
rect 809 113 811 115
rect 805 112 811 113
rect 816 117 820 119
rect 816 115 817 117
rect 819 115 820 117
rect 739 103 762 104
rect 739 101 741 103
rect 743 101 762 103
rect 739 100 762 101
rect 739 94 743 100
rect 698 91 699 93
rect 701 91 702 93
rect 698 86 702 91
rect 698 82 710 86
rect 694 79 695 81
rect 600 68 606 74
rect 706 78 710 82
rect 732 90 743 94
rect 732 84 736 90
rect 758 94 762 100
rect 766 110 770 112
rect 766 108 767 110
rect 769 108 770 110
rect 766 103 770 108
rect 766 101 767 103
rect 769 102 770 103
rect 769 101 782 102
rect 766 98 782 101
rect 778 96 782 98
rect 778 94 783 96
rect 758 93 774 94
rect 758 91 770 93
rect 772 91 774 93
rect 758 90 774 91
rect 778 92 780 94
rect 782 92 783 94
rect 778 90 783 92
rect 732 82 733 84
rect 735 82 736 84
rect 732 80 736 82
rect 778 86 782 90
rect 758 82 782 86
rect 758 79 762 82
rect 706 77 726 78
rect 758 77 759 79
rect 761 77 762 79
rect 706 75 722 77
rect 724 75 726 77
rect 706 74 726 75
rect 745 76 751 77
rect 745 74 747 76
rect 749 74 751 76
rect 758 75 762 77
rect 816 110 820 115
rect 825 117 831 124
rect 855 122 856 124
rect 858 122 859 124
rect 825 115 827 117
rect 829 115 831 117
rect 825 114 831 115
rect 855 117 859 122
rect 911 122 913 124
rect 915 122 917 124
rect 911 121 917 122
rect 855 115 856 117
rect 858 115 859 117
rect 855 113 859 115
rect 863 118 896 119
rect 863 116 892 118
rect 894 116 896 118
rect 863 115 896 116
rect 816 109 817 110
rect 803 108 817 109
rect 819 108 820 110
rect 803 105 820 108
rect 803 93 807 105
rect 863 104 867 115
rect 919 117 936 118
rect 919 115 932 117
rect 934 115 936 117
rect 919 114 936 115
rect 950 115 956 124
rect 844 103 867 104
rect 844 101 846 103
rect 848 101 867 103
rect 844 100 867 101
rect 844 94 848 100
rect 803 91 804 93
rect 806 91 807 93
rect 803 86 807 91
rect 803 82 815 86
rect 799 79 800 81
rect 661 71 667 72
rect 661 69 663 71
rect 665 69 667 71
rect 661 68 667 69
rect 680 71 686 72
rect 680 69 682 71
rect 684 69 686 71
rect 680 68 686 69
rect 745 68 751 74
rect 811 78 815 82
rect 837 90 848 94
rect 837 84 841 90
rect 863 94 867 100
rect 871 110 875 112
rect 871 108 872 110
rect 874 108 875 110
rect 871 103 875 108
rect 871 101 872 103
rect 874 102 875 103
rect 874 101 887 102
rect 871 98 887 101
rect 883 96 887 98
rect 883 94 888 96
rect 863 93 879 94
rect 863 91 875 93
rect 877 91 879 93
rect 863 90 879 91
rect 883 92 885 94
rect 887 92 888 94
rect 883 90 888 92
rect 837 82 838 84
rect 840 82 841 84
rect 837 80 841 82
rect 883 86 887 90
rect 863 82 887 86
rect 863 79 867 82
rect 811 77 831 78
rect 863 77 864 79
rect 866 77 867 79
rect 904 103 905 114
rect 919 110 923 114
rect 950 113 952 115
rect 954 113 956 115
rect 950 112 956 113
rect 961 117 965 119
rect 961 115 962 117
rect 964 115 965 117
rect 908 106 923 110
rect 908 93 912 106
rect 961 110 965 115
rect 970 117 976 124
rect 1000 122 1001 124
rect 1003 122 1004 124
rect 970 115 972 117
rect 974 115 976 117
rect 970 114 976 115
rect 1000 117 1004 122
rect 1000 115 1001 117
rect 1003 115 1004 117
rect 1000 113 1004 115
rect 1008 118 1041 119
rect 1008 116 1037 118
rect 1039 116 1041 118
rect 1008 115 1041 116
rect 1055 115 1061 124
rect 961 109 962 110
rect 948 108 962 109
rect 964 108 965 110
rect 948 105 965 108
rect 927 97 933 98
rect 908 91 909 93
rect 911 91 912 93
rect 908 85 912 91
rect 908 84 926 85
rect 908 82 922 84
rect 924 82 926 84
rect 908 81 926 82
rect 811 75 827 77
rect 829 75 831 77
rect 811 74 831 75
rect 850 76 856 77
rect 850 74 852 76
rect 854 74 856 76
rect 863 75 867 77
rect 948 93 952 105
rect 1008 104 1012 115
rect 1055 113 1057 115
rect 1059 113 1061 115
rect 1055 112 1061 113
rect 1066 117 1070 119
rect 1066 115 1067 117
rect 1069 115 1070 117
rect 989 103 1012 104
rect 989 101 991 103
rect 993 101 1012 103
rect 989 100 1012 101
rect 989 94 993 100
rect 948 91 949 93
rect 951 91 952 93
rect 948 86 952 91
rect 948 82 960 86
rect 944 79 945 81
rect 850 68 856 74
rect 956 78 960 82
rect 982 90 993 94
rect 982 84 986 90
rect 1008 94 1012 100
rect 1016 110 1020 112
rect 1016 108 1017 110
rect 1019 108 1020 110
rect 1016 103 1020 108
rect 1016 101 1017 103
rect 1019 102 1020 103
rect 1019 101 1032 102
rect 1016 98 1032 101
rect 1028 96 1032 98
rect 1028 94 1033 96
rect 1008 93 1024 94
rect 1008 91 1020 93
rect 1022 91 1024 93
rect 1008 90 1024 91
rect 1028 92 1030 94
rect 1032 92 1033 94
rect 1028 90 1033 92
rect 982 82 983 84
rect 985 82 986 84
rect 982 80 986 82
rect 1028 86 1032 90
rect 1008 82 1032 86
rect 1008 79 1012 82
rect 956 77 976 78
rect 1008 77 1009 79
rect 1011 77 1012 79
rect 956 75 972 77
rect 974 75 976 77
rect 956 74 976 75
rect 995 76 1001 77
rect 995 74 997 76
rect 999 74 1001 76
rect 1008 75 1012 77
rect 1066 110 1070 115
rect 1075 117 1081 124
rect 1105 122 1106 124
rect 1108 122 1109 124
rect 1075 115 1077 117
rect 1079 115 1081 117
rect 1075 114 1081 115
rect 1105 117 1109 122
rect 1105 115 1106 117
rect 1108 115 1109 117
rect 1105 113 1109 115
rect 1113 118 1146 119
rect 1113 116 1142 118
rect 1144 116 1146 118
rect 1113 115 1146 116
rect 1066 109 1067 110
rect 1053 108 1067 109
rect 1069 108 1070 110
rect 1053 105 1070 108
rect 1053 93 1057 105
rect 1113 104 1117 115
rect 1094 103 1117 104
rect 1094 101 1096 103
rect 1098 101 1117 103
rect 1094 100 1117 101
rect 1094 94 1098 100
rect 1053 91 1054 93
rect 1056 91 1057 93
rect 1053 86 1057 91
rect 1053 82 1065 86
rect 1049 79 1050 81
rect 911 71 917 72
rect 911 69 913 71
rect 915 69 917 71
rect 911 68 917 69
rect 930 71 936 72
rect 930 69 932 71
rect 934 69 936 71
rect 930 68 936 69
rect 995 68 1001 74
rect 1061 78 1065 82
rect 1087 90 1098 94
rect 1087 84 1091 90
rect 1113 94 1117 100
rect 1121 110 1125 112
rect 1121 108 1122 110
rect 1124 108 1125 110
rect 1121 103 1125 108
rect 1121 101 1122 103
rect 1124 102 1125 103
rect 1124 101 1137 102
rect 1121 98 1137 101
rect 1133 96 1137 98
rect 1133 94 1138 96
rect 1113 93 1129 94
rect 1113 91 1125 93
rect 1127 91 1129 93
rect 1113 90 1129 91
rect 1133 92 1135 94
rect 1137 92 1138 94
rect 1133 90 1138 92
rect 1087 82 1088 84
rect 1090 82 1091 84
rect 1087 80 1091 82
rect 1133 86 1137 90
rect 1113 82 1137 86
rect 1113 79 1117 82
rect 1061 77 1081 78
rect 1113 77 1114 79
rect 1116 77 1117 79
rect 1061 75 1077 77
rect 1079 75 1081 77
rect 1061 74 1081 75
rect 1100 76 1106 77
rect 1100 74 1102 76
rect 1104 74 1106 76
rect 1113 75 1117 77
rect 1100 68 1106 74
rect 160 51 166 52
rect 160 49 162 51
rect 164 49 166 51
rect 160 48 166 49
rect 179 51 185 52
rect 179 49 181 51
rect 183 49 185 51
rect 179 48 185 49
rect 244 46 250 52
rect 205 45 225 46
rect 205 43 221 45
rect 223 43 225 45
rect 244 44 246 46
rect 248 44 250 46
rect 244 43 250 44
rect 257 43 261 45
rect 205 42 225 43
rect 157 38 175 39
rect 157 36 171 38
rect 173 36 175 38
rect 157 35 175 36
rect 157 29 161 35
rect 193 39 194 41
rect 205 38 209 42
rect 257 41 258 43
rect 260 41 261 43
rect 157 27 158 29
rect 160 27 161 29
rect 153 6 154 17
rect 157 14 161 27
rect 176 22 182 23
rect 157 10 172 14
rect 168 6 172 10
rect 197 34 209 38
rect 197 29 201 34
rect 197 27 198 29
rect 200 27 201 29
rect 197 15 201 27
rect 231 38 235 40
rect 231 36 232 38
rect 234 36 235 38
rect 231 30 235 36
rect 257 38 261 41
rect 257 34 281 38
rect 231 26 242 30
rect 238 20 242 26
rect 277 30 281 34
rect 257 29 273 30
rect 257 27 269 29
rect 271 27 273 29
rect 257 26 273 27
rect 277 28 282 30
rect 277 26 279 28
rect 281 26 282 28
rect 257 20 261 26
rect 277 24 282 26
rect 277 22 281 24
rect 238 19 261 20
rect 238 17 240 19
rect 242 17 261 19
rect 238 16 261 17
rect 197 12 214 15
rect 197 11 211 12
rect 210 10 211 11
rect 213 10 214 12
rect 199 7 205 8
rect 168 5 185 6
rect 168 3 181 5
rect 183 3 185 5
rect 168 2 185 3
rect 199 5 201 7
rect 203 5 205 7
rect 160 -2 166 -1
rect 160 -4 162 -2
rect 164 -4 166 -2
rect 199 -4 205 5
rect 210 5 214 10
rect 210 3 211 5
rect 213 3 214 5
rect 210 1 214 3
rect 219 5 225 6
rect 219 3 221 5
rect 223 3 225 5
rect 219 -4 225 3
rect 249 5 253 7
rect 249 3 250 5
rect 252 3 253 5
rect 249 -2 253 3
rect 257 5 261 16
rect 265 19 281 22
rect 265 17 266 19
rect 268 18 281 19
rect 268 17 269 18
rect 265 12 269 17
rect 265 10 266 12
rect 268 10 269 12
rect 265 8 269 10
rect 349 46 355 52
rect 410 51 416 52
rect 410 49 412 51
rect 414 49 416 51
rect 410 48 416 49
rect 429 51 435 52
rect 429 49 431 51
rect 433 49 435 51
rect 429 48 435 49
rect 310 45 330 46
rect 310 43 326 45
rect 328 43 330 45
rect 349 44 351 46
rect 353 44 355 46
rect 349 43 355 44
rect 362 43 366 45
rect 310 42 330 43
rect 298 39 299 41
rect 310 38 314 42
rect 362 41 363 43
rect 365 41 366 43
rect 302 34 314 38
rect 302 29 306 34
rect 302 27 303 29
rect 305 27 306 29
rect 302 15 306 27
rect 336 38 340 40
rect 336 36 337 38
rect 339 36 340 38
rect 336 30 340 36
rect 362 38 366 41
rect 362 34 386 38
rect 336 26 347 30
rect 343 20 347 26
rect 382 30 386 34
rect 362 29 378 30
rect 362 27 374 29
rect 376 27 378 29
rect 362 26 378 27
rect 382 28 387 30
rect 382 26 384 28
rect 386 26 387 28
rect 362 20 366 26
rect 382 24 387 26
rect 382 22 386 24
rect 343 19 366 20
rect 343 17 345 19
rect 347 17 366 19
rect 343 16 366 17
rect 302 12 319 15
rect 302 11 316 12
rect 315 10 316 11
rect 318 10 319 12
rect 304 7 310 8
rect 304 5 306 7
rect 308 5 310 7
rect 257 4 290 5
rect 257 2 286 4
rect 288 2 290 4
rect 257 1 290 2
rect 249 -4 250 -2
rect 252 -4 253 -2
rect 304 -4 310 5
rect 315 5 319 10
rect 315 3 316 5
rect 318 3 319 5
rect 315 1 319 3
rect 324 5 330 6
rect 324 3 326 5
rect 328 3 330 5
rect 324 -4 330 3
rect 354 5 358 7
rect 354 3 355 5
rect 357 3 358 5
rect 354 -2 358 3
rect 362 5 366 16
rect 370 19 386 22
rect 370 17 371 19
rect 373 18 386 19
rect 373 17 374 18
rect 370 12 374 17
rect 494 46 500 52
rect 455 45 475 46
rect 455 43 471 45
rect 473 43 475 45
rect 494 44 496 46
rect 498 44 500 46
rect 494 43 500 44
rect 507 43 511 45
rect 455 42 475 43
rect 370 10 371 12
rect 373 10 374 12
rect 370 8 374 10
rect 407 38 425 39
rect 407 36 421 38
rect 423 36 425 38
rect 407 35 425 36
rect 407 29 411 35
rect 443 39 444 41
rect 455 38 459 42
rect 507 41 508 43
rect 510 41 511 43
rect 407 27 408 29
rect 410 27 411 29
rect 403 6 404 17
rect 407 14 411 27
rect 426 22 432 23
rect 407 10 422 14
rect 418 6 422 10
rect 447 34 459 38
rect 447 29 451 34
rect 447 27 448 29
rect 450 27 451 29
rect 447 15 451 27
rect 481 38 485 40
rect 481 36 482 38
rect 484 36 485 38
rect 481 30 485 36
rect 507 38 511 41
rect 507 34 531 38
rect 481 26 492 30
rect 488 20 492 26
rect 527 30 531 34
rect 507 29 523 30
rect 507 27 519 29
rect 521 27 523 29
rect 507 26 523 27
rect 527 28 532 30
rect 527 26 529 28
rect 531 26 532 28
rect 507 20 511 26
rect 527 24 532 26
rect 527 22 531 24
rect 488 19 511 20
rect 488 17 490 19
rect 492 17 511 19
rect 488 16 511 17
rect 447 12 464 15
rect 447 11 461 12
rect 460 10 461 11
rect 463 10 464 12
rect 449 7 455 8
rect 362 4 395 5
rect 362 2 391 4
rect 393 2 395 4
rect 362 1 395 2
rect 418 5 435 6
rect 418 3 431 5
rect 433 3 435 5
rect 418 2 435 3
rect 449 5 451 7
rect 453 5 455 7
rect 354 -4 355 -2
rect 357 -4 358 -2
rect 410 -2 416 -1
rect 410 -4 412 -2
rect 414 -4 416 -2
rect 449 -4 455 5
rect 460 5 464 10
rect 460 3 461 5
rect 463 3 464 5
rect 460 1 464 3
rect 469 5 475 6
rect 469 3 471 5
rect 473 3 475 5
rect 469 -4 475 3
rect 499 5 503 7
rect 499 3 500 5
rect 502 3 503 5
rect 499 -2 503 3
rect 507 5 511 16
rect 515 19 531 22
rect 515 17 516 19
rect 518 18 531 19
rect 518 17 519 18
rect 515 12 519 17
rect 515 10 516 12
rect 518 10 519 12
rect 515 8 519 10
rect 599 46 605 52
rect 660 51 666 52
rect 660 49 662 51
rect 664 49 666 51
rect 660 48 666 49
rect 679 51 685 52
rect 679 49 681 51
rect 683 49 685 51
rect 679 48 685 49
rect 560 45 580 46
rect 560 43 576 45
rect 578 43 580 45
rect 599 44 601 46
rect 603 44 605 46
rect 599 43 605 44
rect 612 43 616 45
rect 560 42 580 43
rect 548 39 549 41
rect 560 38 564 42
rect 612 41 613 43
rect 615 41 616 43
rect 552 34 564 38
rect 552 29 556 34
rect 552 27 553 29
rect 555 27 556 29
rect 552 15 556 27
rect 586 38 590 40
rect 586 36 587 38
rect 589 36 590 38
rect 586 30 590 36
rect 612 38 616 41
rect 612 34 636 38
rect 586 26 597 30
rect 593 20 597 26
rect 632 30 636 34
rect 612 29 628 30
rect 612 27 624 29
rect 626 27 628 29
rect 612 26 628 27
rect 632 28 637 30
rect 632 26 634 28
rect 636 26 637 28
rect 612 20 616 26
rect 632 24 637 26
rect 632 22 636 24
rect 593 19 616 20
rect 593 17 595 19
rect 597 17 616 19
rect 593 16 616 17
rect 552 12 569 15
rect 552 11 566 12
rect 565 10 566 11
rect 568 10 569 12
rect 554 7 560 8
rect 554 5 556 7
rect 558 5 560 7
rect 507 4 540 5
rect 507 2 536 4
rect 538 2 540 4
rect 507 1 540 2
rect 499 -4 500 -2
rect 502 -4 503 -2
rect 554 -4 560 5
rect 565 5 569 10
rect 565 3 566 5
rect 568 3 569 5
rect 565 1 569 3
rect 574 5 580 6
rect 574 3 576 5
rect 578 3 580 5
rect 574 -4 580 3
rect 604 5 608 7
rect 604 3 605 5
rect 607 3 608 5
rect 604 -2 608 3
rect 612 5 616 16
rect 620 19 636 22
rect 620 17 621 19
rect 623 18 636 19
rect 623 17 624 18
rect 620 12 624 17
rect 744 46 750 52
rect 705 45 725 46
rect 705 43 721 45
rect 723 43 725 45
rect 744 44 746 46
rect 748 44 750 46
rect 744 43 750 44
rect 757 43 761 45
rect 705 42 725 43
rect 620 10 621 12
rect 623 10 624 12
rect 620 8 624 10
rect 657 38 675 39
rect 657 36 671 38
rect 673 36 675 38
rect 657 35 675 36
rect 657 29 661 35
rect 693 39 694 41
rect 705 38 709 42
rect 757 41 758 43
rect 760 41 761 43
rect 657 27 658 29
rect 660 27 661 29
rect 653 6 654 17
rect 657 14 661 27
rect 676 22 682 23
rect 657 10 672 14
rect 668 6 672 10
rect 697 34 709 38
rect 697 29 701 34
rect 697 27 698 29
rect 700 27 701 29
rect 697 15 701 27
rect 731 38 735 40
rect 731 36 732 38
rect 734 36 735 38
rect 731 30 735 36
rect 757 38 761 41
rect 757 34 781 38
rect 731 26 742 30
rect 738 20 742 26
rect 777 30 781 34
rect 757 29 773 30
rect 757 27 769 29
rect 771 27 773 29
rect 757 26 773 27
rect 777 28 782 30
rect 777 26 779 28
rect 781 26 782 28
rect 757 20 761 26
rect 777 24 782 26
rect 777 22 781 24
rect 738 19 761 20
rect 738 17 740 19
rect 742 17 761 19
rect 738 16 761 17
rect 697 12 714 15
rect 697 11 711 12
rect 710 10 711 11
rect 713 10 714 12
rect 699 7 705 8
rect 612 4 645 5
rect 612 2 641 4
rect 643 2 645 4
rect 612 1 645 2
rect 668 5 685 6
rect 668 3 681 5
rect 683 3 685 5
rect 668 2 685 3
rect 699 5 701 7
rect 703 5 705 7
rect 604 -4 605 -2
rect 607 -4 608 -2
rect 660 -2 666 -1
rect 660 -4 662 -2
rect 664 -4 666 -2
rect 699 -4 705 5
rect 710 5 714 10
rect 710 3 711 5
rect 713 3 714 5
rect 710 1 714 3
rect 719 5 725 6
rect 719 3 721 5
rect 723 3 725 5
rect 719 -4 725 3
rect 749 5 753 7
rect 749 3 750 5
rect 752 3 753 5
rect 749 -2 753 3
rect 757 5 761 16
rect 765 19 781 22
rect 765 17 766 19
rect 768 18 781 19
rect 768 17 769 18
rect 765 12 769 17
rect 765 10 766 12
rect 768 10 769 12
rect 765 8 769 10
rect 849 46 855 52
rect 910 51 916 52
rect 910 49 912 51
rect 914 49 916 51
rect 910 48 916 49
rect 929 51 935 52
rect 929 49 931 51
rect 933 49 935 51
rect 929 48 935 49
rect 810 45 830 46
rect 810 43 826 45
rect 828 43 830 45
rect 849 44 851 46
rect 853 44 855 46
rect 849 43 855 44
rect 862 43 866 45
rect 810 42 830 43
rect 798 39 799 41
rect 810 38 814 42
rect 862 41 863 43
rect 865 41 866 43
rect 802 34 814 38
rect 802 29 806 34
rect 802 27 803 29
rect 805 27 806 29
rect 802 15 806 27
rect 836 38 840 40
rect 836 36 837 38
rect 839 36 840 38
rect 836 30 840 36
rect 862 38 866 41
rect 862 34 886 38
rect 836 26 847 30
rect 843 20 847 26
rect 882 30 886 34
rect 862 29 878 30
rect 862 27 874 29
rect 876 27 878 29
rect 862 26 878 27
rect 882 28 887 30
rect 882 26 884 28
rect 886 26 887 28
rect 862 20 866 26
rect 882 24 887 26
rect 882 22 886 24
rect 843 19 866 20
rect 843 17 845 19
rect 847 17 866 19
rect 843 16 866 17
rect 802 12 819 15
rect 802 11 816 12
rect 815 10 816 11
rect 818 10 819 12
rect 804 7 810 8
rect 804 5 806 7
rect 808 5 810 7
rect 757 4 790 5
rect 757 2 786 4
rect 788 2 790 4
rect 757 1 790 2
rect 749 -4 750 -2
rect 752 -4 753 -2
rect 804 -4 810 5
rect 815 5 819 10
rect 815 3 816 5
rect 818 3 819 5
rect 815 1 819 3
rect 824 5 830 6
rect 824 3 826 5
rect 828 3 830 5
rect 824 -4 830 3
rect 854 5 858 7
rect 854 3 855 5
rect 857 3 858 5
rect 854 -2 858 3
rect 862 5 866 16
rect 870 19 886 22
rect 870 17 871 19
rect 873 18 886 19
rect 873 17 874 18
rect 870 12 874 17
rect 994 46 1000 52
rect 955 45 975 46
rect 955 43 971 45
rect 973 43 975 45
rect 994 44 996 46
rect 998 44 1000 46
rect 994 43 1000 44
rect 1007 43 1011 45
rect 955 42 975 43
rect 870 10 871 12
rect 873 10 874 12
rect 870 8 874 10
rect 907 38 925 39
rect 907 36 921 38
rect 923 36 925 38
rect 907 35 925 36
rect 907 29 911 35
rect 943 39 944 41
rect 955 38 959 42
rect 1007 41 1008 43
rect 1010 41 1011 43
rect 907 27 908 29
rect 910 27 911 29
rect 903 6 904 17
rect 907 14 911 27
rect 926 22 932 23
rect 907 10 922 14
rect 918 6 922 10
rect 947 34 959 38
rect 947 29 951 34
rect 947 27 948 29
rect 950 27 951 29
rect 947 15 951 27
rect 981 38 985 40
rect 981 36 982 38
rect 984 36 985 38
rect 981 30 985 36
rect 1007 38 1011 41
rect 1007 34 1031 38
rect 981 26 992 30
rect 988 20 992 26
rect 1027 30 1031 34
rect 1007 29 1023 30
rect 1007 27 1019 29
rect 1021 27 1023 29
rect 1007 26 1023 27
rect 1027 28 1032 30
rect 1027 26 1029 28
rect 1031 26 1032 28
rect 1007 20 1011 26
rect 1027 24 1032 26
rect 1027 22 1031 24
rect 988 19 1011 20
rect 988 17 990 19
rect 992 17 1011 19
rect 988 16 1011 17
rect 947 12 964 15
rect 947 11 961 12
rect 960 10 961 11
rect 963 10 964 12
rect 949 7 955 8
rect 862 4 895 5
rect 862 2 891 4
rect 893 2 895 4
rect 862 1 895 2
rect 918 5 935 6
rect 918 3 931 5
rect 933 3 935 5
rect 918 2 935 3
rect 949 5 951 7
rect 953 5 955 7
rect 854 -4 855 -2
rect 857 -4 858 -2
rect 910 -2 916 -1
rect 910 -4 912 -2
rect 914 -4 916 -2
rect 949 -4 955 5
rect 960 5 964 10
rect 960 3 961 5
rect 963 3 964 5
rect 960 1 964 3
rect 969 5 975 6
rect 969 3 971 5
rect 973 3 975 5
rect 969 -4 975 3
rect 999 5 1003 7
rect 999 3 1000 5
rect 1002 3 1003 5
rect 999 -2 1003 3
rect 1007 5 1011 16
rect 1015 19 1031 22
rect 1015 17 1016 19
rect 1018 18 1031 19
rect 1018 17 1019 18
rect 1015 12 1019 17
rect 1015 10 1016 12
rect 1018 10 1019 12
rect 1015 8 1019 10
rect 1099 46 1105 52
rect 1060 45 1080 46
rect 1060 43 1076 45
rect 1078 43 1080 45
rect 1099 44 1101 46
rect 1103 44 1105 46
rect 1099 43 1105 44
rect 1112 43 1116 45
rect 1060 42 1080 43
rect 1048 39 1049 41
rect 1060 38 1064 42
rect 1112 41 1113 43
rect 1115 41 1116 43
rect 1052 34 1064 38
rect 1052 29 1056 34
rect 1052 27 1053 29
rect 1055 27 1056 29
rect 1052 15 1056 27
rect 1086 38 1090 40
rect 1086 36 1087 38
rect 1089 36 1090 38
rect 1086 30 1090 36
rect 1112 38 1116 41
rect 1112 34 1136 38
rect 1086 26 1097 30
rect 1093 20 1097 26
rect 1132 30 1136 34
rect 1112 29 1128 30
rect 1112 27 1124 29
rect 1126 27 1128 29
rect 1112 26 1128 27
rect 1132 28 1137 30
rect 1132 26 1134 28
rect 1136 26 1137 28
rect 1112 20 1116 26
rect 1132 24 1137 26
rect 1132 22 1136 24
rect 1093 19 1116 20
rect 1093 17 1095 19
rect 1097 17 1116 19
rect 1093 16 1116 17
rect 1052 12 1069 15
rect 1052 11 1066 12
rect 1065 10 1066 11
rect 1068 10 1069 12
rect 1054 7 1060 8
rect 1054 5 1056 7
rect 1058 5 1060 7
rect 1007 4 1040 5
rect 1007 2 1036 4
rect 1038 2 1040 4
rect 1007 1 1040 2
rect 999 -4 1000 -2
rect 1002 -4 1003 -2
rect 1054 -4 1060 5
rect 1065 5 1069 10
rect 1065 3 1066 5
rect 1068 3 1069 5
rect 1065 1 1069 3
rect 1074 5 1080 6
rect 1074 3 1076 5
rect 1078 3 1080 5
rect 1074 -4 1080 3
rect 1104 5 1108 7
rect 1104 3 1105 5
rect 1107 3 1108 5
rect 1104 -2 1108 3
rect 1112 5 1116 16
rect 1120 19 1136 22
rect 1120 17 1121 19
rect 1123 18 1136 19
rect 1123 17 1124 18
rect 1120 12 1124 17
rect 1120 10 1121 12
rect 1123 10 1124 12
rect 1120 8 1124 10
rect 1112 4 1145 5
rect 1112 2 1141 4
rect 1143 2 1145 4
rect 1112 1 1145 2
rect 1104 -4 1105 -2
rect 1107 -4 1108 -2
<< via1 >>
rect 219 315 221 317
rect 234 324 236 326
rect 259 315 261 317
rect 202 299 204 301
rect 242 300 244 302
rect 273 301 275 303
rect 335 324 337 326
rect 362 324 364 326
rect 435 315 437 317
rect 386 312 388 314
rect 354 301 356 303
rect 450 324 452 326
rect 475 315 477 317
rect 418 299 420 301
rect 458 300 460 302
rect 489 301 491 303
rect 551 324 553 326
rect 578 324 580 326
rect 640 315 642 317
rect 602 312 604 314
rect 570 301 572 303
rect 655 324 657 326
rect 680 315 682 317
rect 623 299 625 301
rect 663 300 665 302
rect 694 301 696 303
rect 756 324 758 326
rect 783 324 785 326
rect 859 315 861 317
rect 807 312 809 314
rect 775 301 777 303
rect 874 324 876 326
rect 899 315 901 317
rect 842 299 844 301
rect 882 300 884 302
rect 913 301 915 303
rect 975 324 977 326
rect 1002 324 1004 326
rect 1026 312 1028 314
rect 994 301 996 303
rect 234 252 236 254
rect 242 243 244 245
rect 217 235 219 237
rect 259 235 261 237
rect 274 226 276 228
rect 330 259 332 261
rect 306 226 308 228
rect 333 226 335 228
rect 450 252 452 254
rect 458 243 460 245
rect 433 235 435 237
rect 475 235 477 237
rect 490 226 492 228
rect 546 259 548 261
rect 522 226 524 228
rect 549 226 551 228
rect 655 252 657 254
rect 663 243 665 245
rect 638 235 640 237
rect 680 235 682 237
rect 695 226 697 228
rect 751 259 753 261
rect 727 226 729 228
rect 754 226 756 228
rect 874 252 876 254
rect 882 243 884 245
rect 857 235 859 237
rect 899 235 901 237
rect 914 226 916 228
rect 970 259 972 261
rect 946 226 948 228
rect 973 226 975 228
rect 1070 226 1072 228
rect 1097 226 1099 228
rect 184 154 186 156
rect 216 180 218 182
rect 243 180 245 182
rect 289 180 291 182
rect 321 180 323 182
rect 298 154 300 156
rect 348 180 350 182
rect 331 162 333 164
rect 402 162 404 164
rect 434 154 436 156
rect 466 180 468 182
rect 493 180 495 182
rect 539 180 541 182
rect 571 180 573 182
rect 548 154 550 156
rect 598 180 600 182
rect 583 162 585 164
rect 652 162 654 164
rect 684 154 686 156
rect 716 180 718 182
rect 743 180 745 182
rect 789 180 791 182
rect 821 180 823 182
rect 798 154 800 156
rect 848 180 850 182
rect 833 162 835 164
rect 902 162 904 164
rect 934 154 936 156
rect 966 180 968 182
rect 993 180 995 182
rect 1039 180 1041 182
rect 1071 180 1073 182
rect 1048 154 1050 156
rect 1098 180 1100 182
rect 183 108 185 110
rect 215 82 217 84
rect 242 82 244 84
rect 288 82 290 84
rect 297 108 299 110
rect 330 100 332 102
rect 320 82 322 84
rect 347 82 349 84
rect 433 108 435 110
rect 401 100 403 102
rect 465 82 467 84
rect 492 82 494 84
rect 538 82 540 84
rect 547 108 549 110
rect 582 100 584 102
rect 570 82 572 84
rect 597 82 599 84
rect 683 108 685 110
rect 651 100 653 102
rect 715 82 717 84
rect 742 82 744 84
rect 788 82 790 84
rect 797 108 799 110
rect 832 100 834 102
rect 820 82 822 84
rect 847 82 849 84
rect 933 108 935 110
rect 901 100 903 102
rect 965 82 967 84
rect 992 82 994 84
rect 1038 82 1040 84
rect 1047 108 1049 110
rect 1082 99 1084 101
rect 1070 82 1072 84
rect 1097 82 1099 84
rect 243 64 245 66
rect 493 65 495 67
rect 1082 64 1084 66
rect 492 53 494 55
rect 1081 54 1083 56
rect 182 10 184 12
rect 214 36 216 38
rect 241 36 243 38
rect 287 36 289 38
rect 319 36 321 38
rect 296 10 298 12
rect 346 36 348 38
rect 329 18 331 20
rect 400 18 402 20
rect 432 10 434 12
rect 464 36 466 38
rect 491 36 493 38
rect 537 36 539 38
rect 569 36 571 38
rect 546 10 548 12
rect 596 36 598 38
rect 581 18 583 20
rect 650 18 652 20
rect 682 10 684 12
rect 714 36 716 38
rect 741 36 743 38
rect 787 36 789 38
rect 819 36 821 38
rect 796 10 798 12
rect 846 36 848 38
rect 831 18 833 20
rect 900 18 902 20
rect 932 10 934 12
rect 964 36 966 38
rect 991 36 993 38
rect 1037 36 1039 38
rect 1069 36 1071 38
rect 1046 10 1048 12
rect 1096 36 1098 38
rect 1081 19 1083 21
<< via2 >>
rect 1082 90 1084 92
rect 1082 74 1084 76
rect 1081 44 1083 46
rect 1081 28 1083 30
<< labels >>
rlabel alu1 539 272 539 272 1 Vdd
rlabel alu1 515 272 515 272 6 vdd
rlabel alu1 537 207 537 207 1 Vss
rlabel alu1 435 208 435 208 6 vss
rlabel alu1 435 272 435 272 6 vdd
rlabel alu1 475 208 475 208 4 vss
rlabel alu1 475 272 475 272 4 vdd
rlabel alu1 565 345 565 345 5 Vss
rlabel alu1 587 280 587 280 2 vdd
rlabel alu1 563 280 563 280 5 Vdd
rlabel alu1 435 280 435 280 2 vdd
rlabel alu1 435 344 435 344 2 vss
rlabel alu1 475 344 475 344 2 vss
rlabel alu1 475 280 475 280 2 vdd
rlabel alu1 632 322 632 322 1 a0
rlabel alu1 672 320 672 320 1 a1
rlabel alu1 680 280 680 280 2 vdd
rlabel alu1 680 344 680 344 2 vss
rlabel alu1 640 344 640 344 2 vss
rlabel alu1 640 280 640 280 2 vdd
rlabel alu1 768 280 768 280 5 Vdd
rlabel alu1 792 280 792 280 2 vdd
rlabel alu1 770 345 770 345 5 Vss
rlabel alu1 680 272 680 272 4 vdd
rlabel alu1 680 208 680 208 4 vss
rlabel alu1 672 231 672 231 1 a1
rlabel alu1 648 230 648 230 1 a0
rlabel alu1 640 272 640 272 6 vdd
rlabel alu1 640 208 640 208 6 vss
rlabel alu1 742 207 742 207 1 Vss
rlabel alu1 720 272 720 272 6 vdd
rlabel alu1 744 272 744 272 1 Vdd
rlabel alu1 704 234 704 234 1 p13
rlabel alu1 624 236 624 236 1 p10
rlabel alu1 801 239 801 239 1 p12
rlabel alu1 711 313 711 313 1 p11
rlabel alu1 419 236 419 236 1 p20
rlabel alu1 499 234 499 234 1 p23
rlabel alu1 596 239 596 239 1 p22
rlabel alu1 233 136 233 136 5 Vdd
rlabel alu1 209 136 209 136 8 vdd
rlabel alu1 231 201 231 201 5 Vss
rlabel alu1 338 136 338 136 5 Vdd
rlabel alu1 314 136 314 136 8 vdd
rlabel alu1 336 201 336 201 5 Vss
rlabel alu1 169 136 169 136 8 vdd
rlabel alu1 483 136 483 136 5 Vdd
rlabel alu1 459 136 459 136 8 vdd
rlabel alu1 481 201 481 201 5 Vss
rlabel alu1 588 136 588 136 5 Vdd
rlabel alu1 564 136 564 136 8 vdd
rlabel alu1 586 201 586 201 5 Vss
rlabel alu1 419 136 419 136 8 vdd
rlabel alu1 669 136 669 136 8 vdd
rlabel alu1 836 201 836 201 5 Vss
rlabel alu1 814 136 814 136 8 vdd
rlabel alu1 838 136 838 136 5 Vdd
rlabel alu1 731 201 731 201 5 Vss
rlabel alu1 709 136 709 136 8 vdd
rlabel alu1 733 136 733 136 5 Vdd
rlabel alu1 983 136 983 136 5 Vdd
rlabel alu1 959 136 959 136 8 vdd
rlabel alu1 981 201 981 201 5 Vss
rlabel alu1 1088 136 1088 136 5 Vdd
rlabel alu1 1064 136 1064 136 8 vdd
rlabel alu1 1086 201 1086 201 5 Vss
rlabel alu1 919 136 919 136 8 vdd
rlabel alu1 242 148 242 148 5 p23
rlabel alu1 251 173 251 173 5 p13
rlabel alu1 492 148 492 148 5 p22
rlabel alu1 501 173 501 173 5 p12
rlabel alu1 742 148 742 148 5 p21
rlabel alu1 751 173 751 173 5 p11
rlabel alu1 992 148 992 148 5 p20
rlabel alu1 1001 173 1001 173 5 p10
rlabel via1 656 252 656 252 1 b2
rlabel alu1 664 252 664 252 1 b3
rlabel alu1 672 308 672 308 1 b2
rlabel via1 624 300 624 300 1 b3
rlabel via1 419 300 419 300 1 b1
rlabel alu1 467 308 467 308 1 b0
rlabel via1 451 252 451 252 1 b0
rlabel alu1 459 252 459 252 1 b1
rlabel alu1 443 230 443 230 1 a2
rlabel alu1 467 231 467 231 1 a3
rlabel alu1 427 322 427 322 1 a2
rlabel alu1 467 320 467 320 1 a3
rlabel alu1 506 313 506 313 1 p21
rlabel alu1 1080 156 1080 156 1 Vss
rlabel alu1 153 165 153 165 1 c0
rlabel alu1 395 169 395 169 1 s03
rlabel alu1 645 169 645 169 1 s02
rlabel alu1 895 169 895 169 1 s01
rlabel alu1 1145 169 1145 169 1 s00
rlabel alu1 923 234 923 234 1 p03
rlabel alu1 1020 239 1020 239 1 p02
rlabel alu1 930 313 930 313 1 r1
rlabel alu1 843 236 843 236 1 r0
rlabel via1 843 300 843 300 1 b1
rlabel alu1 851 322 851 322 1 a0
rlabel alu1 891 320 891 320 1 a1
rlabel alu1 891 308 891 308 1 b0
rlabel alu1 899 280 899 280 2 vdd
rlabel alu1 899 344 899 344 2 vss
rlabel alu1 859 344 859 344 2 vss
rlabel alu1 859 280 859 280 2 vdd
rlabel alu1 987 280 987 280 5 Vdd
rlabel alu1 1011 280 1011 280 2 vdd
rlabel alu1 989 345 989 345 5 Vss
rlabel alu1 899 272 899 272 4 vdd
rlabel alu1 899 208 899 208 4 vss
rlabel alu1 891 231 891 231 1 a1
rlabel alu1 883 252 883 252 1 b1
rlabel alu1 875 252 875 252 1 b0
rlabel alu1 867 230 867 230 1 a0
rlabel alu1 859 272 859 272 6 vdd
rlabel alu1 859 208 859 208 6 vss
rlabel alu1 961 207 961 207 1 Vss
rlabel alu1 939 272 939 272 6 vdd
rlabel alu1 963 272 963 272 1 Vdd
rlabel alu1 290 313 290 313 1 p31
rlabel alu1 380 239 380 239 1 p32
rlabel alu1 283 234 283 234 1 p33
rlabel alu1 203 236 203 236 1 p30
rlabel alu1 211 322 211 322 1 a2
rlabel via1 203 300 203 300 1 b3
rlabel alu1 251 320 251 320 1 a3
rlabel alu1 251 308 251 308 1 b2
rlabel alu1 251 231 251 231 1 a3
rlabel alu1 243 252 243 252 1 b3
rlabel via1 235 252 235 252 1 b2
rlabel alu1 227 230 227 230 1 a2
rlabel alu1 259 280 259 280 2 vdd
rlabel alu1 259 344 259 344 2 vss
rlabel alu1 219 344 219 344 2 vss
rlabel alu1 219 280 219 280 2 vdd
rlabel alu1 347 280 347 280 5 Vdd
rlabel alu1 371 280 371 280 2 vdd
rlabel alu1 349 345 349 345 5 Vss
rlabel alu1 259 272 259 272 4 vdd
rlabel alu1 259 208 259 208 4 vss
rlabel alu1 219 272 219 272 6 vdd
rlabel alu1 219 208 219 208 6 vss
rlabel alu1 321 207 321 207 1 Vss
rlabel alu1 299 272 299 272 6 vdd
rlabel alu1 323 272 323 272 1 Vdd
rlabel alu1 232 128 232 128 1 Vdd
rlabel alu1 208 128 208 128 6 vdd
rlabel alu1 230 63 230 63 1 Vss
rlabel alu1 337 128 337 128 1 Vdd
rlabel alu1 313 128 313 128 6 vdd
rlabel alu1 335 63 335 63 1 Vss
rlabel alu1 168 128 168 128 6 vdd
rlabel alu1 482 128 482 128 1 Vdd
rlabel alu1 458 128 458 128 6 vdd
rlabel alu1 480 63 480 63 1 Vss
rlabel alu1 587 128 587 128 1 Vdd
rlabel alu1 563 128 563 128 6 vdd
rlabel alu1 585 63 585 63 1 Vss
rlabel alu1 418 128 418 128 6 vdd
rlabel alu1 668 128 668 128 6 vdd
rlabel alu1 835 63 835 63 1 Vss
rlabel alu1 813 128 813 128 6 vdd
rlabel alu1 837 128 837 128 1 Vdd
rlabel alu1 730 63 730 63 1 Vss
rlabel alu1 708 128 708 128 6 vdd
rlabel alu1 732 128 732 128 1 Vdd
rlabel alu1 982 128 982 128 1 Vdd
rlabel alu1 958 128 958 128 6 vdd
rlabel alu1 980 63 980 63 1 Vss
rlabel alu1 1087 128 1087 128 1 Vdd
rlabel alu1 1063 128 1063 128 6 vdd
rlabel alu1 1085 63 1085 63 1 Vss
rlabel alu1 918 128 918 128 6 vdd
rlabel alu1 1000 91 1000 91 1 p02
rlabel alu1 991 116 991 116 1 s00
rlabel alu1 750 91 750 91 1 p03
rlabel alu1 741 116 741 116 1 s01
rlabel alu1 500 91 500 91 1 Vss
rlabel alu1 491 116 491 116 1 s02
rlabel alu1 250 91 250 91 1 Vss
rlabel alu1 241 116 241 116 1 s03
rlabel alu1 152 99 152 99 1 c1
rlabel alu1 394 95 394 95 1 s13
rlabel alu1 644 95 644 95 1 s12
rlabel alu1 1079 108 1079 108 1 Vss
rlabel alu1 231 -8 231 -8 5 Vdd
rlabel alu1 207 -8 207 -8 8 vdd
rlabel alu1 229 57 229 57 5 Vss
rlabel alu1 336 -8 336 -8 5 Vdd
rlabel alu1 312 -8 312 -8 8 vdd
rlabel alu1 334 57 334 57 5 Vss
rlabel alu1 167 -8 167 -8 8 vdd
rlabel alu1 481 -8 481 -8 5 Vdd
rlabel alu1 457 -8 457 -8 8 vdd
rlabel alu1 479 57 479 57 5 Vss
rlabel alu1 586 -8 586 -8 5 Vdd
rlabel alu1 562 -8 562 -8 8 vdd
rlabel alu1 584 57 584 57 5 Vss
rlabel alu1 417 -8 417 -8 8 vdd
rlabel alu1 667 -8 667 -8 8 vdd
rlabel alu1 834 57 834 57 5 Vss
rlabel alu1 812 -8 812 -8 8 vdd
rlabel alu1 836 -8 836 -8 5 Vdd
rlabel alu1 729 57 729 57 5 Vss
rlabel alu1 707 -8 707 -8 8 vdd
rlabel alu1 731 -8 731 -8 5 Vdd
rlabel alu1 981 -8 981 -8 5 Vdd
rlabel alu1 957 -8 957 -8 8 vdd
rlabel alu1 979 57 979 57 5 Vss
rlabel alu1 1086 -8 1086 -8 5 Vdd
rlabel alu1 1062 -8 1062 -8 8 vdd
rlabel alu1 1084 57 1084 57 5 Vss
rlabel alu1 917 -8 917 -8 8 vdd
rlabel alu1 1078 12 1078 12 5 Vss
rlabel alu1 151 21 151 21 5 c2
rlabel alu1 240 4 240 4 5 p33
rlabel alu1 490 4 490 4 5 p32
rlabel alu1 740 4 740 4 5 p31
rlabel alu1 749 29 749 29 5 s13
rlabel alu1 990 4 990 4 5 p30
rlabel alu1 999 29 999 29 5 s12
rlabel alu1 1143 25 1143 25 5 r4
rlabel alu1 893 25 893 25 5 r5
rlabel alu1 643 25 643 25 5 r6
rlabel alu1 393 25 393 25 5 r7
rlabel alu1 1144 95 1144 95 1 r2
rlabel alu1 894 95 894 95 1 r3
rlabel alu1 1087 272 1087 272 1 Vdd
rlabel alu1 1063 272 1063 272 6 vdd
rlabel alu1 1085 207 1085 207 1 Vss
rlabel alu1 1071 232 1071 232 1 c0
rlabel alu1 1105 235 1105 235 1 c0
rlabel alu1 1096 260 1096 260 1 c1
rlabel alu1 1079 252 1079 252 1 c1
rlabel alu1 249 29 249 29 1 c11
rlabel alu1 1047 234 1047 234 1 c11
rlabel alu1 499 29 499 29 1 sum
rlabel alu1 1144 239 1144 239 1 sum
<< end >>
