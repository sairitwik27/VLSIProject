magic
tech scmos
timestamp 1607599002
<< ab >>
rect 4 54 68 77
rect 6 13 68 54
rect 4 5 68 13
rect 2 0 70 5
rect 2 -8 22 0
rect 3 -72 22 -64
rect 24 -72 64 0
rect 66 -8 70 0
<< nwell >>
rect -1 37 73 82
rect -1 -77 73 -32
<< pwell >>
rect -1 -32 73 37
<< poly >>
rect 21 71 23 75
rect 6 46 12 48
rect 6 44 8 46
rect 10 44 12 46
rect 57 71 59 75
rect 37 62 39 66
rect 47 62 49 66
rect 6 42 12 44
rect 10 41 12 42
rect 21 41 23 44
rect 37 41 39 44
rect 10 39 23 41
rect 29 39 39 41
rect 47 40 49 44
rect 57 41 59 44
rect 13 31 15 39
rect 29 35 31 39
rect 22 33 31 35
rect 43 38 49 40
rect 43 36 45 38
rect 47 36 49 38
rect 43 34 49 36
rect 53 39 59 41
rect 53 37 55 39
rect 57 37 59 39
rect 53 35 59 37
rect 22 31 24 33
rect 26 31 31 33
rect 22 29 31 31
rect 47 31 49 34
rect 29 26 31 29
rect 39 26 41 30
rect 47 29 51 31
rect 49 26 51 29
rect 56 26 58 35
rect 13 19 15 22
rect 13 17 18 19
rect 16 9 18 17
rect 29 13 31 17
rect 39 9 41 17
rect 49 9 51 14
rect 56 9 58 14
rect 16 7 41 9
rect 33 -13 35 -8
rect 40 -13 42 -8
rect 53 -15 55 -11
rect 33 -37 35 -24
rect 40 -29 42 -24
rect 53 -29 55 -24
rect 39 -31 45 -29
rect 39 -33 41 -31
rect 43 -33 45 -31
rect 39 -35 45 -33
rect 49 -31 55 -29
rect 49 -33 51 -31
rect 53 -33 55 -31
rect 49 -35 55 -33
rect 29 -39 35 -37
rect 29 -41 31 -39
rect 33 -41 35 -39
rect 29 -43 35 -41
rect 33 -46 35 -43
rect 43 -46 45 -35
rect 53 -39 55 -35
rect 33 -64 35 -59
rect 43 -64 45 -59
rect 53 -61 55 -57
<< ndif >>
rect 6 29 13 31
rect 6 27 8 29
rect 10 27 13 29
rect 6 25 13 27
rect 8 22 13 25
rect 15 26 20 31
rect 15 22 29 26
rect 20 21 29 22
rect 20 19 22 21
rect 24 19 29 21
rect 20 17 29 19
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 17 39 22
rect 41 22 49 26
rect 41 20 44 22
rect 46 20 49 22
rect 41 17 49 20
rect 44 14 49 17
rect 51 14 56 26
rect 58 14 66 26
rect 60 12 66 14
rect 60 10 62 12
rect 64 10 66 12
rect 60 8 66 10
rect 44 -5 51 -3
rect 44 -7 47 -5
rect 49 -7 51 -5
rect 44 -13 51 -7
rect 26 -15 33 -13
rect 26 -17 28 -15
rect 30 -17 33 -15
rect 26 -19 33 -17
rect 28 -24 33 -19
rect 35 -24 40 -13
rect 42 -15 51 -13
rect 42 -24 53 -15
rect 55 -17 62 -15
rect 55 -19 58 -17
rect 60 -19 62 -17
rect 55 -21 62 -19
rect 55 -24 60 -21
<< pdif >>
rect 16 50 21 71
rect 14 48 21 50
rect 14 46 16 48
rect 18 46 21 48
rect 14 44 21 46
rect 23 69 35 71
rect 23 67 26 69
rect 28 67 35 69
rect 23 62 35 67
rect 52 62 57 71
rect 23 60 26 62
rect 28 60 37 62
rect 23 44 37 60
rect 39 55 47 62
rect 39 53 42 55
rect 44 53 47 55
rect 39 48 47 53
rect 39 46 42 48
rect 44 46 47 48
rect 39 44 47 46
rect 49 55 57 62
rect 49 53 52 55
rect 54 53 57 55
rect 49 44 57 53
rect 59 65 64 71
rect 59 63 66 65
rect 59 61 62 63
rect 64 61 66 63
rect 59 59 66 61
rect 59 44 64 59
rect 47 -46 53 -39
rect 26 -55 33 -46
rect 26 -57 28 -55
rect 30 -57 33 -55
rect 26 -59 33 -57
rect 35 -48 43 -46
rect 35 -50 38 -48
rect 40 -50 43 -48
rect 35 -55 43 -50
rect 35 -57 38 -55
rect 40 -57 43 -55
rect 35 -59 43 -57
rect 45 -53 53 -46
rect 45 -55 48 -53
rect 50 -55 53 -53
rect 45 -57 53 -55
rect 55 -41 62 -39
rect 55 -43 58 -41
rect 60 -43 62 -41
rect 55 -48 62 -43
rect 55 -50 58 -48
rect 60 -50 62 -48
rect 55 -52 62 -50
rect 55 -57 60 -52
rect 45 -59 51 -57
<< alu1 >>
rect 2 72 70 77
rect 2 70 42 72
rect 44 70 70 72
rect 2 69 70 70
rect 6 58 18 64
rect 6 52 11 58
rect 6 50 7 52
rect 9 50 11 52
rect 6 46 11 50
rect 6 44 8 46
rect 10 44 11 46
rect 6 42 11 44
rect 22 33 27 40
rect 50 55 66 56
rect 50 53 52 55
rect 54 53 66 55
rect 50 51 66 53
rect 22 32 24 33
rect 14 31 24 32
rect 26 31 27 33
rect 14 29 27 31
rect 14 27 18 29
rect 20 27 27 29
rect 14 26 27 27
rect 62 23 66 51
rect 42 22 66 23
rect 42 20 44 22
rect 46 20 66 22
rect 42 19 66 20
rect 2 12 70 13
rect 2 10 9 12
rect 11 10 62 12
rect 64 10 70 12
rect 2 -5 70 10
rect 2 -7 47 -5
rect 49 -7 57 -5
rect 59 -7 70 -5
rect 2 -8 70 -7
rect 33 -29 38 -21
rect 50 -17 62 -13
rect 50 -19 58 -17
rect 60 -19 62 -17
rect 33 -31 34 -29
rect 36 -30 38 -29
rect 36 -31 47 -30
rect 33 -33 41 -31
rect 43 -33 47 -31
rect 33 -34 47 -33
rect 26 -39 39 -38
rect 26 -41 31 -39
rect 33 -41 39 -39
rect 26 -42 39 -41
rect 26 -43 30 -42
rect 26 -45 27 -43
rect 29 -45 30 -43
rect 58 -39 62 -19
rect 26 -51 30 -45
rect 57 -41 62 -39
rect 57 -43 58 -41
rect 60 -43 62 -41
rect 57 -48 62 -43
rect 57 -50 58 -48
rect 60 -50 62 -48
rect 57 -52 62 -50
rect 3 -65 66 -64
rect 3 -67 57 -65
rect 59 -67 66 -65
rect 3 -72 66 -67
<< alu2 >>
rect 6 52 11 54
rect 6 50 7 52
rect 9 50 11 52
rect 6 -42 11 50
rect 17 29 21 32
rect 17 27 18 29
rect 20 27 21 29
rect 17 -27 21 27
rect 17 -29 38 -27
rect 17 -31 34 -29
rect 36 -31 38 -29
rect 17 -32 38 -31
rect 6 -43 30 -42
rect 6 -45 27 -43
rect 29 -45 30 -43
rect 6 -46 30 -45
<< ptie >>
rect 7 12 13 14
rect 7 10 9 12
rect 11 10 13 12
rect 7 8 13 10
rect 55 -5 61 -3
rect 55 -7 57 -5
rect 59 -7 61 -5
rect 55 -9 61 -7
<< ntie >>
rect 40 72 46 74
rect 40 70 42 72
rect 44 70 46 72
rect 40 68 46 70
rect 55 -65 61 -63
rect 55 -67 57 -65
rect 59 -67 61 -65
rect 55 -69 61 -67
<< nmos >>
rect 13 22 15 31
rect 29 17 31 26
rect 39 17 41 26
rect 49 14 51 26
rect 56 14 58 26
rect 33 -24 35 -13
rect 40 -24 42 -13
rect 53 -24 55 -15
<< pmos >>
rect 21 44 23 71
rect 37 44 39 62
rect 47 44 49 62
rect 57 44 59 71
rect 33 -59 35 -46
rect 43 -59 45 -46
rect 53 -57 55 -39
<< polyct0 >>
rect 45 36 47 38
rect 55 37 57 39
rect 51 -33 53 -31
<< polyct1 >>
rect 8 44 10 46
rect 24 31 26 33
rect 41 -33 43 -31
rect 31 -41 33 -39
<< ndifct0 >>
rect 8 27 10 29
rect 22 19 24 21
rect 34 22 36 24
rect 28 -17 30 -15
<< ndifct1 >>
rect 44 20 46 22
rect 62 10 64 12
rect 47 -7 49 -5
rect 58 -19 60 -17
<< ntiect1 >>
rect 42 70 44 72
rect 57 -67 59 -65
<< ptiect1 >>
rect 9 10 11 12
rect 57 -7 59 -5
<< pdifct0 >>
rect 16 46 18 48
rect 26 67 28 69
rect 26 60 28 62
rect 42 53 44 55
rect 42 46 44 48
rect 62 61 64 63
rect 28 -57 30 -55
rect 38 -50 40 -48
rect 38 -57 40 -55
rect 48 -55 50 -53
<< pdifct1 >>
rect 52 53 54 55
rect 58 -43 60 -41
rect 58 -50 60 -48
<< alu0 >>
rect 25 67 26 69
rect 28 67 29 69
rect 25 62 29 67
rect 25 60 26 62
rect 28 60 29 62
rect 25 58 29 60
rect 33 63 66 64
rect 33 61 62 63
rect 64 61 66 63
rect 33 60 66 61
rect 33 49 37 60
rect 14 48 37 49
rect 14 46 16 48
rect 18 46 37 48
rect 14 45 37 46
rect 14 39 18 45
rect 7 35 18 39
rect 7 29 11 35
rect 33 39 37 45
rect 41 55 45 57
rect 41 53 42 55
rect 44 53 45 55
rect 41 48 45 53
rect 41 46 42 48
rect 44 47 45 48
rect 44 46 57 47
rect 41 43 57 46
rect 53 41 57 43
rect 53 39 58 41
rect 33 38 49 39
rect 33 36 45 38
rect 47 36 49 38
rect 33 35 49 36
rect 53 37 55 39
rect 57 37 58 39
rect 53 35 58 37
rect 7 27 8 29
rect 10 27 11 29
rect 7 25 11 27
rect 53 31 57 35
rect 33 27 57 31
rect 33 24 37 27
rect 33 22 34 24
rect 36 22 37 24
rect 20 21 26 22
rect 20 19 22 21
rect 24 19 26 21
rect 33 20 37 22
rect 20 13 26 19
rect 26 -15 46 -14
rect 26 -17 28 -15
rect 30 -17 46 -15
rect 26 -18 46 -17
rect 42 -22 46 -18
rect 57 -21 58 -19
rect 42 -26 54 -22
rect 50 -31 54 -26
rect 50 -33 51 -31
rect 53 -33 54 -31
rect 50 -45 54 -33
rect 37 -48 54 -45
rect 37 -50 38 -48
rect 40 -49 54 -48
rect 40 -50 41 -49
rect 26 -55 32 -54
rect 26 -57 28 -55
rect 30 -57 32 -55
rect 26 -64 32 -57
rect 37 -55 41 -50
rect 37 -57 38 -55
rect 40 -57 41 -55
rect 37 -59 41 -57
rect 46 -53 52 -52
rect 46 -55 48 -53
rect 50 -55 52 -53
rect 46 -64 52 -55
<< via1 >>
rect 7 50 9 52
rect 18 27 20 29
rect 34 -31 36 -29
rect 27 -45 29 -43
<< labels >>
rlabel alu1 8 53 8 53 6 b
rlabel alu1 24 33 24 33 6 a
rlabel alu1 36 9 36 9 6 vss
rlabel alu1 36 73 36 73 6 vdd
rlabel alu1 64 42 64 42 1 sum
rlabel alu1 28 -48 28 -48 2 b
rlabel alu1 44 -68 44 -68 2 vdd
rlabel alu1 36 -28 36 -28 2 a
rlabel alu1 44 -4 44 -4 2 vss
rlabel alu1 60 -32 60 -32 1 cout
<< end >>
