magic
tech scmos
timestamp 1607669642
<< ab >>
rect -45 5 -5 77
rect -3 69 2 77
rect 4 69 108 77
rect 4 37 44 69
rect 45 37 108 69
rect 4 5 108 37
rect 118 69 222 77
rect 118 37 158 69
rect 159 37 222 69
rect 118 5 222 37
rect 39 0 45 5
rect 153 0 159 5
<< nwell >>
rect -50 37 227 82
<< pwell >>
rect -50 0 227 37
<< poly >>
rect -23 71 -21 75
rect -16 71 -14 75
rect -36 61 -34 66
rect 61 71 63 75
rect 13 62 15 66
rect 23 64 25 69
rect 33 64 35 69
rect -36 40 -34 43
rect -23 40 -21 50
rect -16 47 -14 50
rect -16 45 -10 47
rect -16 43 -14 45
rect -12 43 -10 45
rect -16 41 -10 43
rect -36 38 -30 40
rect -36 36 -34 38
rect -32 36 -30 38
rect -36 34 -30 36
rect -26 38 -20 40
rect -26 36 -24 38
rect -22 36 -20 38
rect -26 34 -20 36
rect -36 31 -34 34
rect -26 31 -24 34
rect -16 31 -14 41
rect 13 40 15 44
rect 23 40 25 51
rect 33 48 35 51
rect 33 46 39 48
rect 33 44 35 46
rect 37 44 39 46
rect 33 42 39 44
rect 46 46 52 48
rect 46 44 48 46
rect 50 44 52 46
rect 97 71 99 75
rect 77 62 79 66
rect 87 62 89 66
rect 175 71 177 75
rect 127 62 129 66
rect 137 64 139 69
rect 147 64 149 69
rect 46 42 52 44
rect 13 38 19 40
rect 13 36 15 38
rect 17 36 19 38
rect 13 34 19 36
rect 23 38 29 40
rect 23 36 25 38
rect 27 36 29 38
rect 23 34 29 36
rect 13 29 15 34
rect 26 29 28 34
rect 33 29 35 42
rect 50 41 52 42
rect 61 41 63 44
rect 77 41 79 44
rect 50 39 63 41
rect 69 39 79 41
rect 87 40 89 44
rect 97 41 99 44
rect 53 31 55 39
rect 69 35 71 39
rect 62 33 71 35
rect 83 38 89 40
rect 83 36 85 38
rect 87 36 89 38
rect 83 34 89 36
rect 93 39 99 41
rect 93 37 95 39
rect 97 37 99 39
rect 93 35 99 37
rect 127 40 129 44
rect 137 40 139 51
rect 147 48 149 51
rect 147 46 153 48
rect 147 44 149 46
rect 151 44 153 46
rect 147 42 153 44
rect 160 46 166 48
rect 160 44 162 46
rect 164 44 166 46
rect 211 71 213 75
rect 191 62 193 66
rect 201 62 203 66
rect 160 42 166 44
rect 127 38 133 40
rect 127 36 129 38
rect 131 36 133 38
rect 62 31 64 33
rect 66 31 71 33
rect -36 17 -34 22
rect -26 20 -24 25
rect -16 20 -14 25
rect 13 16 15 20
rect 62 29 71 31
rect 87 31 89 34
rect 69 26 71 29
rect 79 26 81 30
rect 87 29 91 31
rect 89 26 91 29
rect 96 26 98 35
rect 127 34 133 36
rect 137 38 143 40
rect 137 36 139 38
rect 141 36 143 38
rect 137 34 143 36
rect 127 29 129 34
rect 140 29 142 34
rect 147 29 149 42
rect 164 41 166 42
rect 175 41 177 44
rect 191 41 193 44
rect 164 39 177 41
rect 183 39 193 41
rect 201 40 203 44
rect 211 41 213 44
rect 167 31 169 39
rect 183 35 185 39
rect 176 33 185 35
rect 197 38 203 40
rect 197 36 199 38
rect 201 36 203 38
rect 197 34 203 36
rect 207 39 213 41
rect 207 37 209 39
rect 211 37 213 39
rect 207 35 213 37
rect 176 31 178 33
rect 180 31 185 33
rect 53 19 55 22
rect 26 13 28 18
rect 33 13 35 18
rect 53 17 58 19
rect 56 9 58 17
rect 69 13 71 17
rect 79 9 81 17
rect 127 16 129 20
rect 176 29 185 31
rect 201 31 203 34
rect 183 26 185 29
rect 193 26 195 30
rect 201 29 205 31
rect 203 26 205 29
rect 210 26 212 35
rect 167 19 169 22
rect 89 9 91 14
rect 96 9 98 14
rect 56 7 81 9
rect 140 13 142 18
rect 147 13 149 18
rect 167 17 172 19
rect 170 9 172 17
rect 183 13 185 17
rect 193 9 195 17
rect 203 9 205 14
rect 210 9 212 14
rect 170 7 195 9
<< ndif >>
rect -43 29 -36 31
rect -43 27 -41 29
rect -39 27 -36 29
rect -43 25 -36 27
rect -41 22 -36 25
rect -34 25 -26 31
rect -24 29 -16 31
rect -24 27 -21 29
rect -19 27 -16 29
rect -24 25 -16 27
rect -14 25 -7 31
rect 46 29 53 31
rect 8 26 13 29
rect -34 22 -28 25
rect -32 18 -28 22
rect -12 18 -7 25
rect 6 24 13 26
rect 6 22 8 24
rect 10 22 13 24
rect 6 20 13 22
rect 15 20 26 29
rect -32 16 -26 18
rect -32 14 -30 16
rect -28 14 -26 16
rect -32 12 -26 14
rect -13 16 -7 18
rect 17 18 26 20
rect 28 18 33 29
rect 35 24 40 29
rect 46 27 48 29
rect 50 27 53 29
rect 46 25 53 27
rect 35 22 42 24
rect 48 22 53 25
rect 55 26 60 31
rect 160 29 167 31
rect 122 26 127 29
rect 55 22 69 26
rect 35 20 38 22
rect 40 20 42 22
rect 35 18 42 20
rect 60 21 69 22
rect 60 19 62 21
rect 64 19 69 21
rect -13 14 -11 16
rect -9 14 -7 16
rect -13 12 -7 14
rect 17 12 24 18
rect 60 17 69 19
rect 71 24 79 26
rect 71 22 74 24
rect 76 22 79 24
rect 71 17 79 22
rect 81 22 89 26
rect 81 20 84 22
rect 86 20 89 22
rect 81 17 89 20
rect 17 10 19 12
rect 21 10 24 12
rect 17 8 24 10
rect 84 14 89 17
rect 91 14 96 26
rect 98 14 106 26
rect 120 24 127 26
rect 120 22 122 24
rect 124 22 127 24
rect 120 20 127 22
rect 129 20 140 29
rect 131 18 140 20
rect 142 18 147 29
rect 149 24 154 29
rect 160 27 162 29
rect 164 27 167 29
rect 160 25 167 27
rect 149 22 156 24
rect 162 22 167 25
rect 169 26 174 31
rect 169 22 183 26
rect 149 20 152 22
rect 154 20 156 22
rect 149 18 156 20
rect 174 21 183 22
rect 174 19 176 21
rect 178 19 183 21
rect 100 12 106 14
rect 100 10 102 12
rect 104 10 106 12
rect 100 8 106 10
rect 131 12 138 18
rect 174 17 183 19
rect 185 24 193 26
rect 185 22 188 24
rect 190 22 193 24
rect 185 17 193 22
rect 195 22 203 26
rect 195 20 198 22
rect 200 20 203 22
rect 195 17 203 20
rect 131 10 133 12
rect 135 10 138 12
rect 131 8 138 10
rect 198 14 203 17
rect 205 14 210 26
rect 212 14 220 26
rect 214 12 220 14
rect 214 10 216 12
rect 218 10 220 12
rect 214 8 220 10
<< pdif >>
rect -32 69 -23 71
rect -32 67 -30 69
rect -28 67 -23 69
rect -32 61 -23 67
rect -43 59 -36 61
rect -43 57 -41 59
rect -39 57 -36 59
rect -43 52 -36 57
rect -43 50 -41 52
rect -39 50 -36 52
rect -43 48 -36 50
rect -41 43 -36 48
rect -34 50 -23 61
rect -21 50 -16 71
rect -14 64 -9 71
rect -14 62 -7 64
rect 17 62 23 64
rect -14 60 -11 62
rect -9 60 -7 62
rect -14 58 -7 60
rect -14 50 -9 58
rect 8 57 13 62
rect 6 55 13 57
rect 6 53 8 55
rect 10 53 13 55
rect -34 43 -26 50
rect 6 48 13 53
rect 6 46 8 48
rect 10 46 13 48
rect 6 44 13 46
rect 15 60 23 62
rect 15 58 18 60
rect 20 58 23 60
rect 15 51 23 58
rect 25 62 33 64
rect 25 60 28 62
rect 30 60 33 62
rect 25 55 33 60
rect 25 53 28 55
rect 30 53 33 55
rect 25 51 33 53
rect 35 62 42 64
rect 35 60 38 62
rect 40 60 42 62
rect 35 51 42 60
rect 15 44 21 51
rect 56 50 61 71
rect 54 48 61 50
rect 54 46 56 48
rect 58 46 61 48
rect 54 44 61 46
rect 63 69 75 71
rect 63 67 66 69
rect 68 67 75 69
rect 63 62 75 67
rect 92 62 97 71
rect 63 60 66 62
rect 68 60 77 62
rect 63 44 77 60
rect 79 55 87 62
rect 79 53 82 55
rect 84 53 87 55
rect 79 48 87 53
rect 79 46 82 48
rect 84 46 87 48
rect 79 44 87 46
rect 89 55 97 62
rect 89 53 92 55
rect 94 53 97 55
rect 89 44 97 53
rect 99 65 104 71
rect 99 63 106 65
rect 99 61 102 63
rect 104 61 106 63
rect 131 62 137 64
rect 99 59 106 61
rect 99 44 104 59
rect 122 57 127 62
rect 120 55 127 57
rect 120 53 122 55
rect 124 53 127 55
rect 120 48 127 53
rect 120 46 122 48
rect 124 46 127 48
rect 120 44 127 46
rect 129 60 137 62
rect 129 58 132 60
rect 134 58 137 60
rect 129 51 137 58
rect 139 62 147 64
rect 139 60 142 62
rect 144 60 147 62
rect 139 55 147 60
rect 139 53 142 55
rect 144 53 147 55
rect 139 51 147 53
rect 149 62 156 64
rect 149 60 152 62
rect 154 60 156 62
rect 149 51 156 60
rect 129 44 135 51
rect 170 50 175 71
rect 168 48 175 50
rect 168 46 170 48
rect 172 46 175 48
rect 168 44 175 46
rect 177 69 189 71
rect 177 67 180 69
rect 182 67 189 69
rect 177 62 189 67
rect 206 62 211 71
rect 177 60 180 62
rect 182 60 191 62
rect 177 44 191 60
rect 193 55 201 62
rect 193 53 196 55
rect 198 53 201 55
rect 193 48 201 53
rect 193 46 196 48
rect 198 46 201 48
rect 193 44 201 46
rect 203 55 211 62
rect 203 53 206 55
rect 208 53 211 55
rect 203 44 211 53
rect 213 65 218 71
rect 213 63 220 65
rect 213 61 216 63
rect 218 61 220 63
rect 213 59 220 61
rect 213 44 218 59
<< alu1 >>
rect -47 72 224 77
rect -47 70 -40 72
rect -38 70 9 72
rect 11 70 82 72
rect 84 70 123 72
rect 125 70 196 72
rect 198 70 224 72
rect -47 69 224 70
rect -43 63 -39 64
rect -43 59 -30 63
rect -43 57 -41 59
rect -43 52 -39 57
rect -43 50 -41 52
rect -43 31 -39 50
rect -11 53 -7 56
rect 6 55 11 57
rect 6 53 8 55
rect 10 53 11 55
rect 46 58 58 64
rect -11 49 11 53
rect -11 47 -7 49
rect -28 45 -7 47
rect -28 43 -14 45
rect -12 43 -7 45
rect 6 48 11 49
rect 6 46 8 48
rect 10 46 11 48
rect 6 44 11 46
rect 38 53 42 56
rect 38 51 39 53
rect 41 51 42 53
rect -43 29 -38 31
rect -43 27 -41 29
rect -39 27 -38 29
rect -43 25 -38 27
rect -28 38 -7 39
rect -28 36 -24 38
rect -22 36 -10 38
rect -8 36 -7 38
rect -28 35 -7 36
rect -11 26 -7 35
rect 6 24 10 44
rect 38 47 42 51
rect 29 46 42 47
rect 29 44 35 46
rect 37 44 42 46
rect 29 43 42 44
rect 46 53 51 58
rect 46 51 48 53
rect 50 51 51 53
rect 46 46 51 51
rect 46 44 48 46
rect 50 44 51 46
rect 46 42 51 44
rect 21 38 35 39
rect 21 36 25 38
rect 27 36 35 38
rect 21 35 35 36
rect 6 22 8 24
rect 10 22 18 24
rect 6 18 18 22
rect 30 29 35 35
rect 30 27 31 29
rect 33 27 35 29
rect 30 26 35 27
rect 62 33 67 40
rect 90 55 106 56
rect 90 53 92 55
rect 94 53 106 55
rect 90 51 106 53
rect 62 32 64 33
rect 54 31 64 32
rect 66 31 67 33
rect 54 29 67 31
rect 54 27 56 29
rect 58 27 67 29
rect 54 26 67 27
rect 102 30 106 51
rect 102 28 103 30
rect 105 28 106 30
rect 102 23 106 28
rect 82 22 106 23
rect 82 20 84 22
rect 86 20 106 22
rect 82 19 106 20
rect 120 55 125 57
rect 120 53 122 55
rect 124 53 125 55
rect 160 58 172 64
rect 120 48 125 53
rect 120 46 122 48
rect 124 46 125 48
rect 120 44 125 46
rect 152 53 156 56
rect 152 51 153 53
rect 155 51 156 53
rect 120 38 124 44
rect 120 36 121 38
rect 123 36 124 38
rect 120 24 124 36
rect 152 47 156 51
rect 143 46 156 47
rect 143 44 149 46
rect 151 44 156 46
rect 143 43 156 44
rect 160 53 165 58
rect 160 51 162 53
rect 164 51 165 53
rect 160 46 165 51
rect 160 44 162 46
rect 164 44 165 46
rect 160 42 165 44
rect 135 38 149 39
rect 135 36 139 38
rect 141 36 149 38
rect 135 35 149 36
rect 120 22 122 24
rect 124 22 132 24
rect 120 18 132 22
rect 144 29 149 35
rect 144 27 145 29
rect 147 27 149 29
rect 144 26 149 27
rect 176 33 181 40
rect 204 55 220 56
rect 204 53 206 55
rect 208 53 220 55
rect 204 51 220 53
rect 176 32 178 33
rect 168 31 178 32
rect 180 31 181 33
rect 168 29 181 31
rect 168 27 170 29
rect 172 27 181 29
rect 168 26 181 27
rect 216 23 220 51
rect 196 22 220 23
rect 196 20 198 22
rect 200 20 220 22
rect 196 19 220 20
rect -47 12 224 13
rect -47 10 -40 12
rect -38 10 9 12
rect 11 10 19 12
rect 21 10 49 12
rect 51 10 102 12
rect 104 10 123 12
rect 125 10 133 12
rect 135 10 163 12
rect 165 10 216 12
rect 218 10 224 12
rect -47 5 224 10
<< alu2 >>
rect 38 53 51 54
rect 38 51 39 53
rect 41 51 48 53
rect 50 51 51 53
rect 38 50 51 51
rect 152 53 165 54
rect 152 51 153 53
rect 155 51 162 53
rect 164 51 165 53
rect 152 50 165 51
rect -11 38 124 39
rect -11 36 -10 38
rect -8 36 121 38
rect 123 36 124 38
rect -11 35 124 36
rect 30 29 62 31
rect 30 27 31 29
rect 33 27 56 29
rect 58 27 62 29
rect 30 26 62 27
rect 102 30 176 31
rect 102 28 103 30
rect 105 29 176 30
rect 105 28 145 29
rect 102 27 145 28
rect 147 27 170 29
rect 172 27 176 29
rect 102 26 176 27
<< ptie >>
rect -42 12 -36 14
rect 7 12 13 14
rect -42 10 -40 12
rect -38 10 -36 12
rect -42 8 -36 10
rect 7 10 9 12
rect 11 10 13 12
rect 7 8 13 10
rect 47 12 53 14
rect 47 10 49 12
rect 51 10 53 12
rect 47 8 53 10
rect 121 12 127 14
rect 121 10 123 12
rect 125 10 127 12
rect 121 8 127 10
rect 161 12 167 14
rect 161 10 163 12
rect 165 10 167 12
rect 161 8 167 10
<< ntie >>
rect -42 72 -36 74
rect -42 70 -40 72
rect -38 70 -36 72
rect 7 72 13 74
rect -42 68 -36 70
rect 7 70 9 72
rect 11 70 13 72
rect 80 72 86 74
rect 7 68 13 70
rect 80 70 82 72
rect 84 70 86 72
rect 121 72 127 74
rect 80 68 86 70
rect 121 70 123 72
rect 125 70 127 72
rect 194 72 200 74
rect 121 68 127 70
rect 194 70 196 72
rect 198 70 200 72
rect 194 68 200 70
<< nmos >>
rect -36 22 -34 31
rect -26 25 -24 31
rect -16 25 -14 31
rect 13 20 15 29
rect 26 18 28 29
rect 33 18 35 29
rect 53 22 55 31
rect 69 17 71 26
rect 79 17 81 26
rect 89 14 91 26
rect 96 14 98 26
rect 127 20 129 29
rect 140 18 142 29
rect 147 18 149 29
rect 167 22 169 31
rect 183 17 185 26
rect 193 17 195 26
rect 203 14 205 26
rect 210 14 212 26
<< pmos >>
rect -36 43 -34 61
rect -23 50 -21 71
rect -16 50 -14 71
rect 13 44 15 62
rect 23 51 25 64
rect 33 51 35 64
rect 61 44 63 71
rect 77 44 79 62
rect 87 44 89 62
rect 97 44 99 71
rect 127 44 129 62
rect 137 51 139 64
rect 147 51 149 64
rect 175 44 177 71
rect 191 44 193 62
rect 201 44 203 62
rect 211 44 213 71
<< polyct0 >>
rect -34 36 -32 38
rect 15 36 17 38
rect 85 36 87 38
rect 95 37 97 39
rect 129 36 131 38
rect 199 36 201 38
rect 209 37 211 39
<< polyct1 >>
rect -14 43 -12 45
rect -24 36 -22 38
rect 35 44 37 46
rect 48 44 50 46
rect 25 36 27 38
rect 149 44 151 46
rect 162 44 164 46
rect 64 31 66 33
rect 139 36 141 38
rect 178 31 180 33
<< ndifct0 >>
rect -21 27 -19 29
rect -30 14 -28 16
rect 48 27 50 29
rect 38 20 40 22
rect 62 19 64 21
rect -11 14 -9 16
rect 74 22 76 24
rect 162 27 164 29
rect 152 20 154 22
rect 176 19 178 21
rect 188 22 190 24
<< ndifct1 >>
rect -41 27 -39 29
rect 8 22 10 24
rect 84 20 86 22
rect 19 10 21 12
rect 122 22 124 24
rect 102 10 104 12
rect 198 20 200 22
rect 133 10 135 12
rect 216 10 218 12
<< ntiect1 >>
rect -40 70 -38 72
rect 9 70 11 72
rect 82 70 84 72
rect 123 70 125 72
rect 196 70 198 72
<< ptiect1 >>
rect -40 10 -38 12
rect 9 10 11 12
rect 49 10 51 12
rect 123 10 125 12
rect 163 10 165 12
<< pdifct0 >>
rect -30 67 -28 69
rect -11 60 -9 62
rect 18 58 20 60
rect 28 60 30 62
rect 28 53 30 55
rect 38 60 40 62
rect 56 46 58 48
rect 66 67 68 69
rect 66 60 68 62
rect 82 53 84 55
rect 82 46 84 48
rect 102 61 104 63
rect 132 58 134 60
rect 142 60 144 62
rect 142 53 144 55
rect 152 60 154 62
rect 170 46 172 48
rect 180 67 182 69
rect 180 60 182 62
rect 196 53 198 55
rect 196 46 198 48
rect 216 61 218 63
<< pdifct1 >>
rect -41 57 -39 59
rect -41 50 -39 52
rect 8 53 10 55
rect 8 46 10 48
rect 92 53 94 55
rect 122 53 124 55
rect 122 46 124 48
rect 206 53 208 55
<< alu0 >>
rect -32 67 -30 69
rect -28 67 -26 69
rect -32 66 -26 67
rect -24 62 -7 63
rect -24 60 -11 62
rect -9 60 -7 62
rect -24 59 -7 60
rect 16 60 22 69
rect -39 48 -38 59
rect -24 55 -20 59
rect 16 58 18 60
rect 20 58 22 60
rect 16 57 22 58
rect 27 62 31 64
rect 27 60 28 62
rect 30 60 31 62
rect -35 51 -20 55
rect 27 55 31 60
rect 36 62 42 69
rect 65 67 66 69
rect 68 67 69 69
rect 36 60 38 62
rect 40 60 42 62
rect 36 59 42 60
rect 65 62 69 67
rect 65 60 66 62
rect 68 60 69 62
rect 65 58 69 60
rect 73 63 106 64
rect 73 61 102 63
rect 104 61 106 63
rect 73 60 106 61
rect 130 60 136 69
rect 27 54 28 55
rect -35 38 -31 51
rect 14 53 28 54
rect 30 53 31 55
rect 14 50 31 53
rect -16 42 -10 43
rect -35 36 -34 38
rect -32 36 -31 38
rect -35 30 -31 36
rect -35 29 -17 30
rect -35 27 -21 29
rect -19 27 -17 29
rect -35 26 -17 27
rect 14 38 18 50
rect 73 49 77 60
rect 130 58 132 60
rect 134 58 136 60
rect 130 57 136 58
rect 141 62 145 64
rect 141 60 142 62
rect 144 60 145 62
rect 54 48 77 49
rect 54 46 56 48
rect 58 46 77 48
rect 54 45 77 46
rect 54 39 58 45
rect 14 36 15 38
rect 17 36 18 38
rect 14 31 18 36
rect 14 27 26 31
rect 10 24 11 26
rect 22 23 26 27
rect 47 35 58 39
rect 47 29 51 35
rect 73 39 77 45
rect 81 55 85 57
rect 81 53 82 55
rect 84 53 85 55
rect 81 48 85 53
rect 81 46 82 48
rect 84 47 85 48
rect 84 46 97 47
rect 81 43 97 46
rect 93 41 97 43
rect 93 39 98 41
rect 73 38 89 39
rect 73 36 85 38
rect 87 36 89 38
rect 73 35 89 36
rect 93 37 95 39
rect 97 37 98 39
rect 93 35 98 37
rect 47 27 48 29
rect 50 27 51 29
rect 47 25 51 27
rect 93 31 97 35
rect 73 27 97 31
rect 73 24 77 27
rect 22 22 42 23
rect 73 22 74 24
rect 76 22 77 24
rect 22 20 38 22
rect 40 20 42 22
rect 22 19 42 20
rect 60 21 66 22
rect 60 19 62 21
rect 64 19 66 21
rect 73 20 77 22
rect 141 55 145 60
rect 150 62 156 69
rect 179 67 180 69
rect 182 67 183 69
rect 150 60 152 62
rect 154 60 156 62
rect 150 59 156 60
rect 179 62 183 67
rect 179 60 180 62
rect 182 60 183 62
rect 179 58 183 60
rect 187 63 220 64
rect 187 61 216 63
rect 218 61 220 63
rect 187 60 220 61
rect 141 54 142 55
rect 128 53 142 54
rect 144 53 145 55
rect 128 50 145 53
rect 128 38 132 50
rect 187 49 191 60
rect 168 48 191 49
rect 168 46 170 48
rect 172 46 191 48
rect 168 45 191 46
rect 168 39 172 45
rect 128 36 129 38
rect 131 36 132 38
rect 128 31 132 36
rect 128 27 140 31
rect 124 24 125 26
rect -32 16 -26 17
rect -32 14 -30 16
rect -28 14 -26 16
rect -32 13 -26 14
rect -13 16 -7 17
rect -13 14 -11 16
rect -9 14 -7 16
rect -13 13 -7 14
rect 60 13 66 19
rect 136 23 140 27
rect 161 35 172 39
rect 161 29 165 35
rect 187 39 191 45
rect 195 55 199 57
rect 195 53 196 55
rect 198 53 199 55
rect 195 48 199 53
rect 195 46 196 48
rect 198 47 199 48
rect 198 46 211 47
rect 195 43 211 46
rect 207 41 211 43
rect 207 39 212 41
rect 187 38 203 39
rect 187 36 199 38
rect 201 36 203 38
rect 187 35 203 36
rect 207 37 209 39
rect 211 37 212 39
rect 207 35 212 37
rect 161 27 162 29
rect 164 27 165 29
rect 161 25 165 27
rect 207 31 211 35
rect 187 27 211 31
rect 187 24 191 27
rect 136 22 156 23
rect 187 22 188 24
rect 190 22 191 24
rect 136 20 152 22
rect 154 20 156 22
rect 136 19 156 20
rect 174 21 180 22
rect 174 19 176 21
rect 178 19 180 21
rect 187 20 191 22
rect 174 13 180 19
<< via1 >>
rect 39 51 41 53
rect -10 36 -8 38
rect 48 51 50 53
rect 31 27 33 29
rect 56 27 58 29
rect 103 28 105 30
rect 153 51 155 53
rect 121 36 123 38
rect 162 51 164 53
rect 145 27 147 29
rect 170 27 172 29
<< labels >>
rlabel alu1 76 9 76 9 6 vss
rlabel alu1 76 73 76 73 6 vdd
rlabel alu1 24 73 24 73 6 vdd
rlabel alu1 24 9 24 9 6 vss
rlabel alu1 190 9 190 9 6 vss
rlabel alu1 190 73 190 73 6 vdd
rlabel alu1 218 33 218 33 1 sum
rlabel alu1 138 73 138 73 6 vdd
rlabel alu1 138 9 138 9 6 vss
rlabel alu1 -25 9 -25 9 6 vss
rlabel alu1 -25 73 -25 73 6 vdd
rlabel alu1 24 36 24 36 1 a
rlabel via1 39 51 39 51 1 b
rlabel alu1 104 33 104 33 1 s1
rlabel via1 155 52 155 52 1 cin
rlabel alu1 -41 39 -41 39 1 cout
<< end >>
