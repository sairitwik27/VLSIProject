magic
tech scmos
timestamp 1608910165
<< ab >>
rect 18 142 66 150
rect 27 77 66 142
rect 68 77 104 150
rect 27 14 64 77
rect 18 6 64 14
rect 66 6 104 77
rect 106 142 111 150
rect 106 86 108 142
rect 106 77 111 86
rect 113 77 176 150
rect 178 118 216 150
rect 178 77 225 118
rect 106 6 146 77
rect 148 6 211 77
rect 216 38 225 77
<< nwell >>
rect 9 38 225 118
<< pwell >>
rect 9 118 225 155
rect 9 1 225 38
<< poly >>
rect 35 137 37 142
rect 42 137 44 142
rect 55 135 57 139
rect 75 137 77 142
rect 82 137 84 142
rect 140 146 165 148
rect 123 141 125 146
rect 130 141 132 146
rect 95 135 97 139
rect 140 138 142 146
rect 150 138 152 142
rect 163 138 165 146
rect 163 136 168 138
rect 187 137 189 142
rect 194 137 196 142
rect 166 133 168 136
rect 35 113 37 126
rect 42 121 44 126
rect 55 121 57 126
rect 41 119 47 121
rect 41 117 43 119
rect 45 117 47 119
rect 41 115 47 117
rect 51 119 57 121
rect 51 117 53 119
rect 55 117 57 119
rect 51 115 57 117
rect 31 111 37 113
rect 31 109 33 111
rect 35 109 37 111
rect 31 107 37 109
rect 35 104 37 107
rect 45 104 47 115
rect 55 111 57 115
rect 75 113 77 126
rect 82 121 84 126
rect 95 121 97 126
rect 81 119 87 121
rect 81 117 83 119
rect 85 117 87 119
rect 81 115 87 117
rect 91 119 97 121
rect 123 120 125 129
rect 130 126 132 129
rect 130 124 134 126
rect 140 125 142 129
rect 150 126 152 129
rect 132 121 134 124
rect 150 124 159 126
rect 207 135 209 139
rect 150 122 155 124
rect 157 122 159 124
rect 91 117 93 119
rect 95 117 97 119
rect 91 115 97 117
rect 71 111 77 113
rect 71 109 73 111
rect 75 109 77 111
rect 71 107 77 109
rect 75 104 77 107
rect 85 104 87 115
rect 95 111 97 115
rect 122 118 128 120
rect 122 116 124 118
rect 126 116 128 118
rect 122 114 128 116
rect 132 119 138 121
rect 132 117 134 119
rect 136 117 138 119
rect 132 115 138 117
rect 150 120 159 122
rect 150 116 152 120
rect 166 116 168 124
rect 122 111 124 114
rect 132 111 134 115
rect 142 114 152 116
rect 158 114 171 116
rect 142 111 144 114
rect 158 111 160 114
rect 169 113 171 114
rect 187 113 189 126
rect 194 121 196 126
rect 207 121 209 126
rect 193 119 199 121
rect 193 117 195 119
rect 197 117 199 119
rect 193 115 199 117
rect 203 119 209 121
rect 203 117 205 119
rect 207 117 209 119
rect 203 115 209 117
rect 169 111 175 113
rect 35 86 37 91
rect 45 86 47 91
rect 55 89 57 93
rect 75 86 77 91
rect 85 86 87 91
rect 95 89 97 93
rect 132 89 134 93
rect 142 89 144 93
rect 122 80 124 84
rect 169 109 171 111
rect 173 109 175 111
rect 169 107 175 109
rect 183 111 189 113
rect 183 109 185 111
rect 187 109 189 111
rect 183 107 189 109
rect 187 104 189 107
rect 197 104 199 115
rect 207 111 209 115
rect 187 86 189 91
rect 197 86 199 91
rect 207 89 209 93
rect 158 80 160 84
rect 35 63 37 67
rect 45 65 47 70
rect 55 65 57 70
rect 75 65 77 70
rect 85 65 87 70
rect 164 72 166 76
rect 95 63 97 67
rect 115 63 117 67
rect 125 65 127 70
rect 135 65 137 70
rect 35 41 37 45
rect 45 41 47 52
rect 55 49 57 52
rect 75 49 77 52
rect 55 47 61 49
rect 55 45 57 47
rect 59 45 61 47
rect 55 43 61 45
rect 71 47 77 49
rect 71 45 73 47
rect 75 45 77 47
rect 71 43 77 45
rect 35 39 41 41
rect 35 37 37 39
rect 39 37 41 39
rect 35 35 41 37
rect 45 39 51 41
rect 45 37 47 39
rect 49 37 51 39
rect 45 35 51 37
rect 35 30 37 35
rect 48 30 50 35
rect 55 30 57 43
rect 75 30 77 43
rect 85 41 87 52
rect 95 41 97 45
rect 81 39 87 41
rect 81 37 83 39
rect 85 37 87 39
rect 81 35 87 37
rect 91 39 97 41
rect 91 37 93 39
rect 95 37 97 39
rect 91 35 97 37
rect 82 30 84 35
rect 95 30 97 35
rect 115 41 117 45
rect 125 41 127 52
rect 135 49 137 52
rect 135 47 141 49
rect 135 45 137 47
rect 139 45 141 47
rect 135 43 141 45
rect 149 47 155 49
rect 149 45 151 47
rect 153 45 155 47
rect 200 72 202 76
rect 180 63 182 67
rect 190 63 192 67
rect 149 43 155 45
rect 115 39 121 41
rect 115 37 117 39
rect 119 37 121 39
rect 115 35 121 37
rect 125 39 131 41
rect 125 37 127 39
rect 129 37 131 39
rect 125 35 131 37
rect 115 30 117 35
rect 128 30 130 35
rect 135 30 137 43
rect 153 42 155 43
rect 164 42 166 45
rect 180 42 182 45
rect 153 40 166 42
rect 172 40 182 42
rect 190 41 192 45
rect 200 42 202 45
rect 156 32 158 40
rect 172 36 174 40
rect 165 34 174 36
rect 186 39 192 41
rect 186 37 188 39
rect 190 37 192 39
rect 186 35 192 37
rect 196 40 202 42
rect 196 38 198 40
rect 200 38 202 40
rect 196 36 202 38
rect 165 32 167 34
rect 169 32 174 34
rect 35 17 37 21
rect 48 14 50 19
rect 55 14 57 19
rect 75 14 77 19
rect 82 14 84 19
rect 95 17 97 21
rect 115 17 117 21
rect 165 30 174 32
rect 190 32 192 35
rect 172 27 174 30
rect 182 27 184 31
rect 190 30 194 32
rect 192 27 194 30
rect 199 27 201 36
rect 156 20 158 23
rect 128 14 130 19
rect 135 14 137 19
rect 156 18 161 20
rect 159 10 161 18
rect 172 14 174 18
rect 182 10 184 18
rect 192 10 194 15
rect 199 10 201 15
rect 159 8 184 10
<< ndif >>
rect 46 145 53 147
rect 46 143 49 145
rect 51 143 53 145
rect 46 137 53 143
rect 86 145 93 147
rect 86 143 89 145
rect 91 143 93 145
rect 28 135 35 137
rect 28 133 30 135
rect 32 133 35 135
rect 28 131 35 133
rect 30 126 35 131
rect 37 126 42 137
rect 44 135 53 137
rect 86 137 93 143
rect 115 145 121 147
rect 115 143 117 145
rect 119 143 121 145
rect 115 141 121 143
rect 68 135 75 137
rect 44 126 55 135
rect 57 133 64 135
rect 57 131 60 133
rect 62 131 64 133
rect 68 133 70 135
rect 72 133 75 135
rect 68 131 75 133
rect 57 129 64 131
rect 57 126 62 129
rect 70 126 75 131
rect 77 126 82 137
rect 84 135 93 137
rect 84 126 95 135
rect 97 133 104 135
rect 97 131 100 133
rect 102 131 104 133
rect 97 129 104 131
rect 115 129 123 141
rect 125 129 130 141
rect 132 138 137 141
rect 198 145 205 147
rect 198 143 201 145
rect 203 143 205 145
rect 132 135 140 138
rect 132 133 135 135
rect 137 133 140 135
rect 132 129 140 133
rect 142 133 150 138
rect 142 131 145 133
rect 147 131 150 133
rect 142 129 150 131
rect 152 136 161 138
rect 198 137 205 143
rect 152 134 157 136
rect 159 134 161 136
rect 152 133 161 134
rect 180 135 187 137
rect 180 133 182 135
rect 184 133 187 135
rect 152 129 166 133
rect 97 126 102 129
rect 161 124 166 129
rect 168 130 173 133
rect 180 131 187 133
rect 168 128 175 130
rect 168 126 171 128
rect 173 126 175 128
rect 182 126 187 131
rect 189 126 194 137
rect 196 135 205 137
rect 196 126 207 135
rect 209 133 216 135
rect 209 131 212 133
rect 214 131 216 133
rect 209 129 216 131
rect 209 126 214 129
rect 168 124 175 126
rect 149 30 156 32
rect 30 27 35 30
rect 28 25 35 27
rect 28 23 30 25
rect 32 23 35 25
rect 28 21 35 23
rect 37 21 48 30
rect 39 19 48 21
rect 50 19 55 30
rect 57 25 62 30
rect 70 25 75 30
rect 57 23 64 25
rect 57 21 60 23
rect 62 21 64 23
rect 57 19 64 21
rect 68 23 75 25
rect 68 21 70 23
rect 72 21 75 23
rect 68 19 75 21
rect 77 19 82 30
rect 84 21 95 30
rect 97 27 102 30
rect 110 27 115 30
rect 97 25 104 27
rect 97 23 100 25
rect 102 23 104 25
rect 97 21 104 23
rect 108 25 115 27
rect 108 23 110 25
rect 112 23 115 25
rect 108 21 115 23
rect 117 21 128 30
rect 84 19 93 21
rect 39 13 46 19
rect 39 11 41 13
rect 43 11 46 13
rect 39 9 46 11
rect 86 13 93 19
rect 119 19 128 21
rect 130 19 135 30
rect 137 25 142 30
rect 149 28 151 30
rect 153 28 156 30
rect 149 26 156 28
rect 137 23 144 25
rect 151 23 156 26
rect 158 27 163 32
rect 158 23 172 27
rect 137 21 140 23
rect 142 21 144 23
rect 137 19 144 21
rect 163 22 172 23
rect 163 20 165 22
rect 167 20 172 22
rect 86 11 89 13
rect 91 11 93 13
rect 86 9 93 11
rect 119 13 126 19
rect 163 18 172 20
rect 174 25 182 27
rect 174 23 177 25
rect 179 23 182 25
rect 174 18 182 23
rect 184 23 192 27
rect 184 21 187 23
rect 189 21 192 23
rect 184 18 192 21
rect 119 11 121 13
rect 123 11 126 13
rect 119 9 126 11
rect 187 15 192 18
rect 194 15 199 27
rect 201 15 209 27
rect 203 13 209 15
rect 203 11 205 13
rect 207 11 209 13
rect 203 9 209 11
<< pdif >>
rect 49 104 55 111
rect 28 95 35 104
rect 28 93 30 95
rect 32 93 35 95
rect 28 91 35 93
rect 37 102 45 104
rect 37 100 40 102
rect 42 100 45 102
rect 37 95 45 100
rect 37 93 40 95
rect 42 93 45 95
rect 37 91 45 93
rect 47 97 55 104
rect 47 95 50 97
rect 52 95 55 97
rect 47 93 55 95
rect 57 109 64 111
rect 57 107 60 109
rect 62 107 64 109
rect 57 102 64 107
rect 89 104 95 111
rect 57 100 60 102
rect 62 100 64 102
rect 57 98 64 100
rect 57 93 62 98
rect 68 95 75 104
rect 68 93 70 95
rect 72 93 75 95
rect 47 91 53 93
rect 68 91 75 93
rect 77 102 85 104
rect 77 100 80 102
rect 82 100 85 102
rect 77 95 85 100
rect 77 93 80 95
rect 82 93 85 95
rect 77 91 85 93
rect 87 97 95 104
rect 87 95 90 97
rect 92 95 95 97
rect 87 93 95 95
rect 97 109 104 111
rect 97 107 100 109
rect 102 107 104 109
rect 97 102 104 107
rect 97 100 100 102
rect 102 100 104 102
rect 97 98 104 100
rect 97 93 102 98
rect 117 96 122 111
rect 115 94 122 96
rect 87 91 93 93
rect 115 92 117 94
rect 119 92 122 94
rect 115 90 122 92
rect 117 84 122 90
rect 124 102 132 111
rect 124 100 127 102
rect 129 100 132 102
rect 124 93 132 100
rect 134 109 142 111
rect 134 107 137 109
rect 139 107 142 109
rect 134 102 142 107
rect 134 100 137 102
rect 139 100 142 102
rect 134 93 142 100
rect 144 95 158 111
rect 144 93 153 95
rect 155 93 158 95
rect 124 84 129 93
rect 146 88 158 93
rect 146 86 153 88
rect 155 86 158 88
rect 146 84 158 86
rect 160 109 167 111
rect 160 107 163 109
rect 165 107 167 109
rect 160 105 167 107
rect 160 84 165 105
rect 201 104 207 111
rect 180 95 187 104
rect 180 93 182 95
rect 184 93 187 95
rect 180 91 187 93
rect 189 102 197 104
rect 189 100 192 102
rect 194 100 197 102
rect 189 95 197 100
rect 189 93 192 95
rect 194 93 197 95
rect 189 91 197 93
rect 199 97 207 104
rect 199 95 202 97
rect 204 95 207 97
rect 199 93 207 95
rect 209 109 216 111
rect 209 107 212 109
rect 214 107 216 109
rect 209 102 216 107
rect 209 100 212 102
rect 214 100 216 102
rect 209 98 216 100
rect 209 93 214 98
rect 199 91 205 93
rect 39 63 45 65
rect 30 58 35 63
rect 28 56 35 58
rect 28 54 30 56
rect 32 54 35 56
rect 28 49 35 54
rect 28 47 30 49
rect 32 47 35 49
rect 28 45 35 47
rect 37 61 45 63
rect 37 59 40 61
rect 42 59 45 61
rect 37 52 45 59
rect 47 63 55 65
rect 47 61 50 63
rect 52 61 55 63
rect 47 56 55 61
rect 47 54 50 56
rect 52 54 55 56
rect 47 52 55 54
rect 57 63 64 65
rect 57 61 60 63
rect 62 61 64 63
rect 57 52 64 61
rect 68 63 75 65
rect 68 61 70 63
rect 72 61 75 63
rect 68 52 75 61
rect 77 63 85 65
rect 77 61 80 63
rect 82 61 85 63
rect 77 56 85 61
rect 77 54 80 56
rect 82 54 85 56
rect 77 52 85 54
rect 87 63 93 65
rect 119 63 125 65
rect 87 61 95 63
rect 87 59 90 61
rect 92 59 95 61
rect 87 52 95 59
rect 37 45 43 52
rect 89 45 95 52
rect 97 58 102 63
rect 110 58 115 63
rect 97 56 104 58
rect 97 54 100 56
rect 102 54 104 56
rect 97 49 104 54
rect 97 47 100 49
rect 102 47 104 49
rect 97 45 104 47
rect 108 56 115 58
rect 108 54 110 56
rect 112 54 115 56
rect 108 49 115 54
rect 108 47 110 49
rect 112 47 115 49
rect 108 45 115 47
rect 117 61 125 63
rect 117 59 120 61
rect 122 59 125 61
rect 117 52 125 59
rect 127 63 135 65
rect 127 61 130 63
rect 132 61 135 63
rect 127 56 135 61
rect 127 54 130 56
rect 132 54 135 56
rect 127 52 135 54
rect 137 63 144 65
rect 137 61 140 63
rect 142 61 144 63
rect 137 52 144 61
rect 117 45 123 52
rect 159 51 164 72
rect 157 49 164 51
rect 157 47 159 49
rect 161 47 164 49
rect 157 45 164 47
rect 166 70 178 72
rect 166 68 169 70
rect 171 68 178 70
rect 166 63 178 68
rect 195 63 200 72
rect 166 61 169 63
rect 171 61 180 63
rect 166 45 180 61
rect 182 56 190 63
rect 182 54 185 56
rect 187 54 190 56
rect 182 49 190 54
rect 182 47 185 49
rect 187 47 190 49
rect 182 45 190 47
rect 192 56 200 63
rect 192 54 195 56
rect 197 54 200 56
rect 192 45 200 54
rect 202 66 207 72
rect 202 64 209 66
rect 202 62 205 64
rect 207 62 209 64
rect 202 60 209 62
rect 202 45 207 60
<< alu1 >>
rect 18 145 216 150
rect 18 143 49 145
rect 51 143 59 145
rect 61 143 89 145
rect 91 143 99 145
rect 101 143 117 145
rect 119 143 170 145
rect 172 143 201 145
rect 203 143 211 145
rect 213 143 216 145
rect 18 142 216 143
rect 35 120 40 129
rect 52 133 64 137
rect 52 131 60 133
rect 62 131 64 133
rect 60 128 64 131
rect 35 119 49 120
rect 35 117 43 119
rect 45 117 46 119
rect 48 117 49 119
rect 35 116 49 117
rect 28 111 41 112
rect 28 109 33 111
rect 35 109 41 111
rect 28 108 41 109
rect 28 103 32 108
rect 60 126 61 128
rect 63 126 64 128
rect 60 111 64 126
rect 75 120 80 129
rect 92 133 104 137
rect 92 131 100 133
rect 102 131 104 133
rect 75 119 89 120
rect 75 117 83 119
rect 85 117 86 119
rect 88 117 89 119
rect 75 116 89 117
rect 28 101 29 103
rect 31 101 32 103
rect 28 99 32 101
rect 59 109 64 111
rect 59 107 60 109
rect 62 107 64 109
rect 59 102 64 107
rect 59 100 60 102
rect 62 100 64 102
rect 59 98 64 100
rect 68 111 81 112
rect 68 109 73 111
rect 75 109 81 111
rect 68 108 81 109
rect 68 104 72 108
rect 100 111 104 131
rect 68 102 69 104
rect 71 102 72 104
rect 68 99 72 102
rect 99 109 104 111
rect 99 107 100 109
rect 102 107 104 109
rect 99 105 104 107
rect 99 103 100 105
rect 102 103 104 105
rect 99 102 104 103
rect 99 100 100 102
rect 102 100 104 102
rect 99 98 104 100
rect 115 135 139 136
rect 115 133 135 135
rect 137 133 139 135
rect 115 132 139 133
rect 115 104 119 132
rect 154 128 167 129
rect 154 126 162 128
rect 164 126 167 128
rect 154 124 167 126
rect 154 122 155 124
rect 157 123 167 124
rect 157 122 159 123
rect 115 102 131 104
rect 115 100 127 102
rect 129 100 131 102
rect 115 99 131 100
rect 154 115 159 122
rect 187 128 192 129
rect 187 126 189 128
rect 191 126 192 128
rect 187 120 192 126
rect 204 133 216 137
rect 204 131 212 133
rect 214 131 216 133
rect 187 119 201 120
rect 187 117 195 119
rect 197 117 201 119
rect 187 116 201 117
rect 170 112 175 113
rect 170 111 176 112
rect 180 111 193 112
rect 170 109 171 111
rect 173 109 185 111
rect 187 109 193 111
rect 170 108 193 109
rect 170 106 184 108
rect 170 97 175 106
rect 180 105 184 106
rect 212 116 216 131
rect 212 114 213 116
rect 215 114 216 116
rect 212 111 216 114
rect 180 103 181 105
rect 183 103 184 105
rect 180 99 184 103
rect 211 109 216 111
rect 211 107 212 109
rect 214 107 216 109
rect 211 102 216 107
rect 163 91 175 97
rect 211 100 212 102
rect 214 100 216 102
rect 211 98 216 100
rect 27 85 216 86
rect 27 83 59 85
rect 61 83 99 85
rect 101 83 137 85
rect 139 83 211 85
rect 213 83 216 85
rect 27 73 216 83
rect 27 71 31 73
rect 33 71 99 73
rect 101 71 111 73
rect 113 71 185 73
rect 187 71 216 73
rect 27 70 216 71
rect 28 56 33 58
rect 28 54 30 56
rect 32 54 33 56
rect 28 49 33 54
rect 28 47 30 49
rect 32 47 33 49
rect 28 45 33 47
rect 60 56 64 57
rect 60 54 61 56
rect 63 54 64 56
rect 28 25 32 45
rect 60 48 64 54
rect 51 47 64 48
rect 51 45 57 47
rect 59 45 64 47
rect 51 44 64 45
rect 68 48 72 57
rect 99 56 104 58
rect 68 47 81 48
rect 68 45 69 47
rect 71 45 73 47
rect 75 45 81 47
rect 68 44 81 45
rect 43 39 57 40
rect 43 37 44 39
rect 46 37 47 39
rect 49 37 57 39
rect 43 36 57 37
rect 28 23 30 25
rect 32 23 40 25
rect 28 19 40 23
rect 52 27 57 36
rect 75 39 89 40
rect 75 37 83 39
rect 85 37 86 39
rect 88 37 89 39
rect 75 36 89 37
rect 99 54 100 56
rect 102 54 104 56
rect 99 49 104 54
rect 99 47 100 49
rect 102 47 104 49
rect 99 45 104 47
rect 75 27 80 36
rect 100 30 104 45
rect 100 28 101 30
rect 103 28 104 30
rect 100 25 104 28
rect 92 23 100 25
rect 102 23 104 25
rect 92 19 104 23
rect 108 56 113 58
rect 108 54 110 56
rect 112 54 113 56
rect 149 63 161 65
rect 149 61 157 63
rect 159 61 161 63
rect 149 59 161 61
rect 108 49 113 54
rect 108 47 110 49
rect 112 47 113 49
rect 108 45 113 47
rect 108 25 112 45
rect 140 50 144 57
rect 149 50 154 59
rect 140 48 154 50
rect 131 47 154 48
rect 131 45 137 47
rect 139 45 151 47
rect 153 45 154 47
rect 131 44 144 45
rect 148 44 154 45
rect 149 43 154 44
rect 123 39 137 40
rect 123 37 127 39
rect 129 37 137 39
rect 123 36 137 37
rect 108 23 110 25
rect 112 23 120 25
rect 108 19 120 23
rect 132 30 137 36
rect 132 28 133 30
rect 135 28 137 30
rect 132 27 137 28
rect 165 34 170 41
rect 193 56 209 57
rect 193 54 195 56
rect 197 54 209 56
rect 193 52 209 54
rect 165 33 167 34
rect 157 32 167 33
rect 169 32 170 34
rect 157 30 170 32
rect 157 28 160 30
rect 162 28 170 30
rect 157 27 170 28
rect 205 24 209 52
rect 185 23 209 24
rect 185 21 187 23
rect 189 21 209 23
rect 185 20 209 21
rect 18 13 213 14
rect 18 11 31 13
rect 33 11 41 13
rect 43 11 89 13
rect 91 11 99 13
rect 101 11 111 13
rect 113 11 121 13
rect 123 11 152 13
rect 154 11 205 13
rect 207 11 213 13
rect 18 6 213 11
<< alu2 >>
rect 60 128 192 129
rect 60 126 61 128
rect 63 126 162 128
rect 164 126 189 128
rect 191 126 192 128
rect 60 125 192 126
rect 43 119 49 120
rect 43 117 46 119
rect 48 117 49 119
rect 20 103 32 104
rect 20 101 29 103
rect 31 101 32 103
rect 20 99 32 101
rect 20 26 25 99
rect 43 39 49 117
rect 85 119 89 120
rect 85 117 86 119
rect 88 117 89 119
rect 68 104 72 105
rect 68 102 69 104
rect 71 102 72 104
rect 68 78 72 102
rect 60 74 72 78
rect 60 56 64 74
rect 60 54 61 56
rect 63 54 64 56
rect 60 53 64 54
rect 43 37 44 39
rect 46 37 49 39
rect 43 36 49 37
rect 68 47 72 48
rect 68 45 69 47
rect 71 45 72 47
rect 68 26 72 45
rect 85 39 89 117
rect 212 116 216 120
rect 212 114 213 116
rect 215 114 216 116
rect 99 105 184 106
rect 99 103 100 105
rect 102 103 181 105
rect 183 103 184 105
rect 99 102 184 103
rect 212 79 216 114
rect 156 74 216 79
rect 156 63 161 74
rect 156 61 157 63
rect 159 61 161 63
rect 156 59 161 61
rect 85 37 86 39
rect 88 37 89 39
rect 85 36 89 37
rect 100 30 165 31
rect 100 28 101 30
rect 103 28 133 30
rect 135 28 160 30
rect 162 28 165 30
rect 100 27 165 28
rect 100 26 138 27
rect 20 22 72 26
<< ptie >>
rect 57 145 63 147
rect 57 143 59 145
rect 61 143 63 145
rect 57 141 63 143
rect 97 145 103 147
rect 97 143 99 145
rect 101 143 103 145
rect 97 141 103 143
rect 168 145 174 147
rect 168 143 170 145
rect 172 143 174 145
rect 168 141 174 143
rect 209 145 215 147
rect 209 143 211 145
rect 213 143 215 145
rect 209 141 215 143
rect 29 13 35 15
rect 29 11 31 13
rect 33 11 35 13
rect 29 9 35 11
rect 97 13 103 15
rect 97 11 99 13
rect 101 11 103 13
rect 97 9 103 11
rect 109 13 115 15
rect 109 11 111 13
rect 113 11 115 13
rect 109 9 115 11
rect 150 13 156 15
rect 150 11 152 13
rect 154 11 156 13
rect 150 9 156 11
<< ntie >>
rect 57 85 63 87
rect 57 83 59 85
rect 61 83 63 85
rect 57 81 63 83
rect 97 85 103 87
rect 97 83 99 85
rect 101 83 103 85
rect 135 85 141 87
rect 97 81 103 83
rect 135 83 137 85
rect 139 83 141 85
rect 209 85 215 87
rect 135 81 141 83
rect 209 83 211 85
rect 213 83 215 85
rect 209 81 215 83
rect 29 73 35 75
rect 29 71 31 73
rect 33 71 35 73
rect 29 69 35 71
rect 97 73 103 75
rect 97 71 99 73
rect 101 71 103 73
rect 97 69 103 71
rect 109 73 115 75
rect 109 71 111 73
rect 113 71 115 73
rect 183 73 189 75
rect 109 69 115 71
rect 183 71 185 73
rect 187 71 189 73
rect 183 69 189 71
<< nmos >>
rect 35 126 37 137
rect 42 126 44 137
rect 55 126 57 135
rect 75 126 77 137
rect 82 126 84 137
rect 95 126 97 135
rect 123 129 125 141
rect 130 129 132 141
rect 140 129 142 138
rect 150 129 152 138
rect 166 124 168 133
rect 187 126 189 137
rect 194 126 196 137
rect 207 126 209 135
rect 35 21 37 30
rect 48 19 50 30
rect 55 19 57 30
rect 75 19 77 30
rect 82 19 84 30
rect 95 21 97 30
rect 115 21 117 30
rect 128 19 130 30
rect 135 19 137 30
rect 156 23 158 32
rect 172 18 174 27
rect 182 18 184 27
rect 192 15 194 27
rect 199 15 201 27
<< pmos >>
rect 35 91 37 104
rect 45 91 47 104
rect 55 93 57 111
rect 75 91 77 104
rect 85 91 87 104
rect 95 93 97 111
rect 122 84 124 111
rect 132 93 134 111
rect 142 93 144 111
rect 158 84 160 111
rect 187 91 189 104
rect 197 91 199 104
rect 207 93 209 111
rect 35 45 37 63
rect 45 52 47 65
rect 55 52 57 65
rect 75 52 77 65
rect 85 52 87 65
rect 95 45 97 63
rect 115 45 117 63
rect 125 52 127 65
rect 135 52 137 65
rect 164 45 166 72
rect 180 45 182 63
rect 190 45 192 63
rect 200 45 202 72
<< polyct0 >>
rect 53 117 55 119
rect 93 117 95 119
rect 124 116 126 118
rect 134 117 136 119
rect 205 117 207 119
rect 37 37 39 39
rect 93 37 95 39
rect 117 37 119 39
rect 188 37 190 39
rect 198 38 200 40
<< polyct1 >>
rect 43 117 45 119
rect 33 109 35 111
rect 83 117 85 119
rect 155 122 157 124
rect 73 109 75 111
rect 195 117 197 119
rect 171 109 173 111
rect 185 109 187 111
rect 57 45 59 47
rect 73 45 75 47
rect 47 37 49 39
rect 83 37 85 39
rect 137 45 139 47
rect 151 45 153 47
rect 127 37 129 39
rect 167 32 169 34
<< ndifct0 >>
rect 30 133 32 135
rect 70 133 72 135
rect 145 131 147 133
rect 157 134 159 136
rect 182 133 184 135
rect 171 126 173 128
rect 60 21 62 23
rect 70 21 72 23
rect 151 28 153 30
rect 140 21 142 23
rect 165 20 167 22
rect 177 23 179 25
<< ndifct1 >>
rect 49 143 51 145
rect 89 143 91 145
rect 117 143 119 145
rect 60 131 62 133
rect 100 131 102 133
rect 201 143 203 145
rect 135 133 137 135
rect 212 131 214 133
rect 30 23 32 25
rect 100 23 102 25
rect 110 23 112 25
rect 41 11 43 13
rect 89 11 91 13
rect 187 21 189 23
rect 121 11 123 13
rect 205 11 207 13
<< ntiect1 >>
rect 59 83 61 85
rect 99 83 101 85
rect 137 83 139 85
rect 211 83 213 85
rect 31 71 33 73
rect 99 71 101 73
rect 111 71 113 73
rect 185 71 187 73
<< ptiect1 >>
rect 59 143 61 145
rect 99 143 101 145
rect 170 143 172 145
rect 211 143 213 145
rect 31 11 33 13
rect 99 11 101 13
rect 111 11 113 13
rect 152 11 154 13
<< pdifct0 >>
rect 30 93 32 95
rect 40 100 42 102
rect 40 93 42 95
rect 50 95 52 97
rect 70 93 72 95
rect 80 100 82 102
rect 80 93 82 95
rect 90 95 92 97
rect 117 92 119 94
rect 137 107 139 109
rect 137 100 139 102
rect 153 93 155 95
rect 153 86 155 88
rect 163 107 165 109
rect 182 93 184 95
rect 192 100 194 102
rect 192 93 194 95
rect 202 95 204 97
rect 40 59 42 61
rect 50 61 52 63
rect 50 54 52 56
rect 60 61 62 63
rect 70 61 72 63
rect 80 61 82 63
rect 80 54 82 56
rect 90 59 92 61
rect 120 59 122 61
rect 130 61 132 63
rect 130 54 132 56
rect 140 61 142 63
rect 159 47 161 49
rect 169 68 171 70
rect 169 61 171 63
rect 185 54 187 56
rect 185 47 187 49
rect 205 62 207 64
<< pdifct1 >>
rect 60 107 62 109
rect 60 100 62 102
rect 100 107 102 109
rect 100 100 102 102
rect 127 100 129 102
rect 212 107 214 109
rect 212 100 214 102
rect 30 54 32 56
rect 30 47 32 49
rect 100 54 102 56
rect 100 47 102 49
rect 110 54 112 56
rect 110 47 112 49
rect 195 54 197 56
<< alu0 >>
rect 28 135 48 136
rect 28 133 30 135
rect 32 133 48 135
rect 28 132 48 133
rect 44 128 48 132
rect 68 135 88 136
rect 68 133 70 135
rect 72 133 88 135
rect 68 132 88 133
rect 59 129 60 131
rect 44 124 56 128
rect 52 119 56 124
rect 52 117 53 119
rect 55 117 56 119
rect 52 105 56 117
rect 84 128 88 132
rect 155 136 161 142
rect 99 129 100 131
rect 84 124 96 128
rect 92 119 96 124
rect 92 117 93 119
rect 95 117 96 119
rect 39 102 56 105
rect 39 100 40 102
rect 42 101 56 102
rect 42 100 43 101
rect 28 95 34 96
rect 28 93 30 95
rect 32 93 34 95
rect 28 86 34 93
rect 39 95 43 100
rect 92 105 96 117
rect 79 102 96 105
rect 79 100 80 102
rect 82 101 96 102
rect 82 100 83 101
rect 39 93 40 95
rect 42 93 43 95
rect 39 91 43 93
rect 48 97 54 98
rect 48 95 50 97
rect 52 95 54 97
rect 48 86 54 95
rect 68 95 74 96
rect 68 93 70 95
rect 72 93 74 95
rect 68 86 74 93
rect 79 95 83 100
rect 144 133 148 135
rect 155 134 157 136
rect 159 134 161 136
rect 155 133 161 134
rect 180 135 200 136
rect 180 133 182 135
rect 184 133 200 135
rect 144 131 145 133
rect 147 131 148 133
rect 180 132 200 133
rect 144 128 148 131
rect 124 124 148 128
rect 124 120 128 124
rect 170 128 174 130
rect 170 126 171 128
rect 173 126 174 128
rect 123 118 128 120
rect 123 116 124 118
rect 126 116 128 118
rect 132 119 148 120
rect 132 117 134 119
rect 136 117 148 119
rect 132 116 148 117
rect 123 114 128 116
rect 124 112 128 114
rect 124 109 140 112
rect 124 108 137 109
rect 136 107 137 108
rect 139 107 140 109
rect 136 102 140 107
rect 136 100 137 102
rect 139 100 140 102
rect 136 98 140 100
rect 144 110 148 116
rect 170 120 174 126
rect 163 116 174 120
rect 196 128 200 132
rect 211 129 212 131
rect 196 124 208 128
rect 204 119 208 124
rect 204 117 205 119
rect 207 117 208 119
rect 163 110 167 116
rect 144 109 167 110
rect 144 107 163 109
rect 165 107 167 109
rect 144 106 167 107
rect 79 93 80 95
rect 82 93 83 95
rect 79 91 83 93
rect 88 97 94 98
rect 88 95 90 97
rect 92 95 94 97
rect 144 95 148 106
rect 204 105 208 117
rect 191 102 208 105
rect 191 100 192 102
rect 194 101 208 102
rect 194 100 195 101
rect 88 86 94 95
rect 115 94 148 95
rect 115 92 117 94
rect 119 92 148 94
rect 115 91 148 92
rect 152 95 156 97
rect 152 93 153 95
rect 155 93 156 95
rect 152 88 156 93
rect 180 95 186 96
rect 180 93 182 95
rect 184 93 186 95
rect 152 86 153 88
rect 155 86 156 88
rect 180 86 186 93
rect 191 95 195 100
rect 191 93 192 95
rect 194 93 195 95
rect 191 91 195 93
rect 200 97 206 98
rect 200 95 202 97
rect 204 95 206 97
rect 200 86 206 95
rect 38 61 44 70
rect 38 59 40 61
rect 42 59 44 61
rect 38 58 44 59
rect 49 63 53 65
rect 49 61 50 63
rect 52 61 53 63
rect 49 56 53 61
rect 58 63 64 70
rect 58 61 60 63
rect 62 61 64 63
rect 58 60 64 61
rect 68 63 74 70
rect 68 61 70 63
rect 72 61 74 63
rect 68 60 74 61
rect 79 63 83 65
rect 79 61 80 63
rect 82 61 83 63
rect 49 55 50 56
rect 36 54 50 55
rect 52 54 53 56
rect 36 51 53 54
rect 36 39 40 51
rect 79 56 83 61
rect 88 61 94 70
rect 88 59 90 61
rect 92 59 94 61
rect 88 58 94 59
rect 118 61 124 70
rect 118 59 120 61
rect 122 59 124 61
rect 118 58 124 59
rect 129 63 133 65
rect 129 61 130 63
rect 132 61 133 63
rect 79 54 80 56
rect 82 55 83 56
rect 82 54 96 55
rect 79 51 96 54
rect 36 37 37 39
rect 39 37 40 39
rect 36 32 40 37
rect 36 28 48 32
rect 32 25 33 27
rect 44 24 48 28
rect 92 39 96 51
rect 92 37 93 39
rect 95 37 96 39
rect 92 32 96 37
rect 84 28 96 32
rect 84 24 88 28
rect 99 25 100 27
rect 44 23 64 24
rect 44 21 60 23
rect 62 21 64 23
rect 44 20 64 21
rect 68 23 88 24
rect 68 21 70 23
rect 72 21 88 23
rect 68 20 88 21
rect 129 56 133 61
rect 138 63 144 70
rect 168 68 169 70
rect 171 68 172 70
rect 138 61 140 63
rect 142 61 144 63
rect 138 60 144 61
rect 168 63 172 68
rect 168 61 169 63
rect 171 61 172 63
rect 168 59 172 61
rect 176 64 209 65
rect 176 62 205 64
rect 207 62 209 64
rect 176 61 209 62
rect 129 55 130 56
rect 116 54 130 55
rect 132 54 133 56
rect 116 51 133 54
rect 116 39 120 51
rect 176 50 180 61
rect 157 49 180 50
rect 157 47 159 49
rect 161 47 180 49
rect 157 46 180 47
rect 157 40 161 46
rect 116 37 117 39
rect 119 37 120 39
rect 116 32 120 37
rect 116 28 128 32
rect 112 25 113 27
rect 124 24 128 28
rect 150 36 161 40
rect 150 30 154 36
rect 176 40 180 46
rect 184 56 188 58
rect 184 54 185 56
rect 187 54 188 56
rect 184 49 188 54
rect 184 47 185 49
rect 187 48 188 49
rect 187 47 200 48
rect 184 44 200 47
rect 196 42 200 44
rect 196 40 201 42
rect 176 39 192 40
rect 176 37 188 39
rect 190 37 192 39
rect 176 36 192 37
rect 196 38 198 40
rect 200 38 201 40
rect 196 36 201 38
rect 150 28 151 30
rect 153 28 154 30
rect 150 26 154 28
rect 196 32 200 36
rect 176 28 200 32
rect 176 25 180 28
rect 124 23 144 24
rect 176 23 177 25
rect 179 23 180 25
rect 124 21 140 23
rect 142 21 144 23
rect 124 20 144 21
rect 163 22 169 23
rect 163 20 165 22
rect 167 20 169 22
rect 176 21 180 23
rect 163 14 169 20
<< via1 >>
rect 46 117 48 119
rect 61 126 63 128
rect 86 117 88 119
rect 29 101 31 103
rect 69 102 71 104
rect 100 103 102 105
rect 162 126 164 128
rect 189 126 191 128
rect 213 114 215 116
rect 181 103 183 105
rect 61 54 63 56
rect 69 45 71 47
rect 44 37 46 39
rect 86 37 88 39
rect 101 28 103 30
rect 157 61 159 63
rect 133 28 135 30
rect 160 28 162 30
<< labels >>
rlabel alu1 150 74 150 74 1 Vdd
rlabel alu1 126 74 126 74 6 vdd
rlabel alu1 148 9 148 9 1 Vss
rlabel alu1 46 10 46 10 6 vss
rlabel alu1 46 74 46 74 6 vdd
rlabel alu1 54 32 54 32 1 a0
rlabel alu1 62 54 62 54 1 b0
rlabel alu1 30 38 30 38 1 p0
rlabel alu1 70 54 70 54 1 b1
rlabel alu1 78 33 78 33 1 a1
rlabel alu1 86 10 86 10 4 vss
rlabel alu1 86 74 86 74 4 vdd
rlabel alu1 176 147 176 147 5 Vss
rlabel alu1 198 82 198 82 2 vdd
rlabel alu1 174 82 174 82 5 Vdd
rlabel alu1 207 41 207 41 1 p2
rlabel alu1 117 115 117 115 1 p1
rlabel alu1 110 36 110 36 1 p3
rlabel alu1 46 82 46 82 2 vdd
rlabel alu1 46 146 46 146 2 vss
rlabel alu1 86 146 86 146 2 vss
rlabel alu1 86 82 86 82 2 vdd
rlabel alu1 78 110 78 110 1 b0
rlabel alu1 78 122 78 122 1 a1
rlabel alu1 38 124 38 124 1 a0
rlabel via1 30 102 30 102 1 b1
<< end >>
