magic
tech scmos
timestamp 1607889199
<< ab >>
rect 88 581 94 586
rect 202 581 208 586
rect 4 5 44 581
rect 53 549 157 581
rect 53 517 93 549
rect 94 517 157 549
rect 46 501 51 517
rect 53 501 157 517
rect 53 469 93 501
rect 94 469 157 501
rect 53 405 157 469
rect 53 373 93 405
rect 94 373 157 405
rect 46 357 51 373
rect 53 357 157 373
rect 53 325 93 357
rect 94 325 157 357
rect 53 261 157 325
rect 53 229 93 261
rect 94 229 157 261
rect 46 213 51 229
rect 53 213 157 229
rect 53 181 93 213
rect 94 181 157 213
rect 53 117 157 181
rect 53 85 93 117
rect 94 85 157 117
rect 46 69 51 85
rect 53 69 157 85
rect 53 37 93 69
rect 94 37 157 69
rect 53 5 157 37
rect 167 549 271 581
rect 272 573 276 581
rect 167 517 207 549
rect 208 517 271 549
rect 167 501 271 517
rect 272 501 274 517
rect 167 469 207 501
rect 208 469 271 501
rect 167 405 271 469
rect 272 429 276 445
rect 167 373 207 405
rect 208 373 271 405
rect 167 357 271 373
rect 272 357 274 373
rect 167 325 207 357
rect 208 325 271 357
rect 167 261 271 325
rect 272 285 276 301
rect 167 229 207 261
rect 208 229 271 261
rect 167 213 271 229
rect 272 213 274 229
rect 167 181 207 213
rect 208 181 271 213
rect 167 117 271 181
rect 272 141 276 157
rect 167 85 207 117
rect 208 85 271 117
rect 167 69 271 85
rect 272 69 274 85
rect 167 37 207 69
rect 208 37 271 69
rect 167 5 271 37
rect 272 5 276 13
rect 278 5 318 581
rect 319 573 383 581
rect 322 517 383 573
rect 319 501 383 517
rect 322 445 383 501
rect 319 429 383 445
rect 322 373 383 429
rect 319 357 383 373
rect 322 301 383 357
rect 319 285 383 301
rect 322 229 383 285
rect 319 213 383 229
rect 322 157 383 213
rect 319 141 383 157
rect 322 85 383 141
rect 319 69 383 85
rect 322 13 383 69
rect 319 5 383 13
rect 387 5 451 581
rect 455 5 518 581
rect 520 573 560 581
rect 562 573 632 581
rect 521 517 560 573
rect 563 517 626 573
rect 520 501 560 517
rect 561 501 626 517
rect 627 501 632 517
rect 521 445 560 501
rect 563 445 626 501
rect 520 429 560 445
rect 562 429 632 445
rect 521 373 560 429
rect 563 373 626 429
rect 520 357 560 373
rect 561 357 626 373
rect 627 357 632 373
rect 521 301 560 357
rect 563 301 626 357
rect 520 285 560 301
rect 562 285 632 301
rect 521 229 560 285
rect 563 229 626 285
rect 520 213 560 229
rect 561 213 626 229
rect 627 213 632 229
rect 521 157 560 213
rect 563 157 626 213
rect 520 141 560 157
rect 562 141 632 157
rect 521 85 560 141
rect 563 85 626 141
rect 520 69 560 85
rect 561 69 626 85
rect 627 69 632 85
rect 521 13 560 69
rect 563 13 626 69
rect 520 5 560 13
rect 562 5 632 13
rect 88 0 94 5
rect 202 0 208 5
<< nwell >>
rect -1 469 632 549
rect -1 325 632 405
rect -1 181 632 261
rect -1 37 632 117
<< pwell >>
rect -1 549 632 586
rect -1 405 632 469
rect -1 261 632 325
rect -1 117 632 181
rect -1 0 632 37
<< poly >>
rect 13 564 15 569
rect 23 561 25 566
rect 33 561 35 566
rect 62 566 64 570
rect 75 568 77 573
rect 82 568 84 573
rect 105 577 130 579
rect 105 569 107 577
rect 118 569 120 573
rect 128 569 130 577
rect 138 572 140 577
rect 145 572 147 577
rect 102 567 107 569
rect 102 564 104 567
rect 13 552 15 555
rect 23 552 25 555
rect 13 550 19 552
rect 13 548 15 550
rect 17 548 19 550
rect 13 546 19 548
rect 23 550 29 552
rect 23 548 25 550
rect 27 548 29 550
rect 23 546 29 548
rect 13 543 15 546
rect 26 536 28 546
rect 33 545 35 555
rect 62 552 64 557
rect 75 552 77 557
rect 62 550 68 552
rect 62 548 64 550
rect 66 548 68 550
rect 62 546 68 548
rect 72 550 78 552
rect 72 548 74 550
rect 76 548 78 550
rect 72 546 78 548
rect 33 543 39 545
rect 33 541 35 543
rect 37 541 39 543
rect 62 542 64 546
rect 33 539 39 541
rect 33 536 35 539
rect 13 520 15 525
rect 72 535 74 546
rect 82 544 84 557
rect 176 566 178 570
rect 189 568 191 573
rect 196 568 198 573
rect 219 577 244 579
rect 219 569 221 577
rect 232 569 234 573
rect 242 569 244 577
rect 252 572 254 577
rect 259 572 261 577
rect 118 557 120 560
rect 111 555 120 557
rect 128 556 130 560
rect 138 557 140 560
rect 102 547 104 555
rect 111 553 113 555
rect 115 553 120 555
rect 111 551 120 553
rect 136 555 140 557
rect 136 552 138 555
rect 118 547 120 551
rect 132 550 138 552
rect 145 551 147 560
rect 216 567 221 569
rect 216 564 218 567
rect 176 552 178 557
rect 189 552 191 557
rect 132 548 134 550
rect 136 548 138 550
rect 99 545 112 547
rect 118 545 128 547
rect 132 546 138 548
rect 99 544 101 545
rect 82 542 88 544
rect 82 540 84 542
rect 86 540 88 542
rect 82 538 88 540
rect 95 542 101 544
rect 110 542 112 545
rect 126 542 128 545
rect 136 542 138 546
rect 142 549 148 551
rect 142 547 144 549
rect 146 547 148 549
rect 142 545 148 547
rect 146 542 148 545
rect 176 550 182 552
rect 176 548 178 550
rect 180 548 182 550
rect 176 546 182 548
rect 186 550 192 552
rect 186 548 188 550
rect 190 548 192 550
rect 186 546 192 548
rect 176 542 178 546
rect 95 540 97 542
rect 99 540 101 542
rect 95 538 101 540
rect 82 535 84 538
rect 62 520 64 524
rect 72 517 74 522
rect 82 517 84 522
rect 26 511 28 515
rect 33 511 35 515
rect 126 520 128 524
rect 136 520 138 524
rect 110 511 112 515
rect 186 535 188 546
rect 196 544 198 557
rect 287 568 289 573
rect 294 568 296 573
rect 329 577 348 579
rect 232 557 234 560
rect 225 555 234 557
rect 242 556 244 560
rect 252 557 254 560
rect 216 547 218 555
rect 225 553 227 555
rect 229 553 234 555
rect 225 551 234 553
rect 250 555 254 557
rect 250 552 252 555
rect 232 547 234 551
rect 246 550 252 552
rect 259 551 261 560
rect 307 566 309 570
rect 329 567 331 577
rect 339 569 341 573
rect 346 569 348 577
rect 423 577 442 579
rect 356 569 358 574
rect 363 569 365 574
rect 373 569 375 574
rect 396 569 398 574
rect 406 569 408 574
rect 413 569 415 574
rect 423 569 425 577
rect 430 569 432 573
rect 246 548 248 550
rect 250 548 252 550
rect 213 545 226 547
rect 232 545 242 547
rect 246 546 252 548
rect 213 544 215 545
rect 196 542 202 544
rect 196 540 198 542
rect 200 540 202 542
rect 196 538 202 540
rect 209 542 215 544
rect 224 542 226 545
rect 240 542 242 545
rect 250 542 252 546
rect 256 549 262 551
rect 256 547 258 549
rect 260 547 262 549
rect 256 545 262 547
rect 260 542 262 545
rect 287 544 289 557
rect 294 552 296 557
rect 307 552 309 557
rect 293 550 299 552
rect 293 548 295 550
rect 297 548 299 550
rect 293 546 299 548
rect 303 550 309 552
rect 303 548 305 550
rect 307 548 309 550
rect 303 546 309 548
rect 283 542 289 544
rect 209 540 211 542
rect 213 540 215 542
rect 209 538 215 540
rect 196 535 198 538
rect 176 520 178 524
rect 186 517 188 522
rect 196 517 198 522
rect 146 511 148 515
rect 240 520 242 524
rect 250 520 252 524
rect 224 511 226 515
rect 283 540 285 542
rect 287 540 289 542
rect 283 538 289 540
rect 287 535 289 538
rect 297 535 299 546
rect 307 542 309 546
rect 329 543 331 561
rect 339 552 341 561
rect 335 550 341 552
rect 335 548 337 550
rect 339 548 341 550
rect 335 546 341 548
rect 346 548 348 561
rect 356 558 358 561
rect 352 556 358 558
rect 352 554 354 556
rect 356 554 358 556
rect 352 552 358 554
rect 346 546 358 548
rect 363 547 365 561
rect 440 567 442 577
rect 490 577 509 579
rect 463 569 465 574
rect 473 569 475 574
rect 480 569 482 574
rect 490 569 492 577
rect 497 569 499 573
rect 373 557 375 560
rect 396 557 398 560
rect 370 555 376 557
rect 370 553 372 555
rect 374 553 376 555
rect 370 551 376 553
rect 395 555 401 557
rect 395 553 397 555
rect 399 553 401 555
rect 395 551 401 553
rect 329 532 331 535
rect 322 530 331 532
rect 339 531 341 546
rect 345 540 351 542
rect 345 538 347 540
rect 349 538 351 540
rect 345 536 351 538
rect 346 531 348 536
rect 356 531 358 546
rect 362 545 368 547
rect 362 543 364 545
rect 366 543 368 545
rect 362 541 368 543
rect 363 531 365 541
rect 373 533 375 551
rect 396 533 398 551
rect 406 547 408 561
rect 413 558 415 561
rect 413 556 419 558
rect 413 554 415 556
rect 417 554 419 556
rect 413 552 419 554
rect 423 548 425 561
rect 403 545 409 547
rect 403 543 405 545
rect 407 543 409 545
rect 403 541 409 543
rect 413 546 425 548
rect 430 552 432 561
rect 430 550 436 552
rect 430 548 432 550
rect 434 548 436 550
rect 430 546 436 548
rect 322 528 324 530
rect 326 528 328 530
rect 322 526 328 528
rect 287 517 289 522
rect 297 517 299 522
rect 307 520 309 524
rect 260 511 262 515
rect 406 531 408 541
rect 413 531 415 546
rect 420 540 426 542
rect 420 538 422 540
rect 424 538 426 540
rect 420 536 426 538
rect 423 531 425 536
rect 430 531 432 546
rect 440 543 442 561
rect 507 567 509 577
rect 589 577 614 579
rect 529 564 531 569
rect 463 557 465 560
rect 462 555 468 557
rect 462 553 464 555
rect 466 553 468 555
rect 462 551 468 553
rect 440 532 442 535
rect 463 533 465 551
rect 473 547 475 561
rect 480 558 482 561
rect 480 556 486 558
rect 480 554 482 556
rect 484 554 486 556
rect 480 552 486 554
rect 490 548 492 561
rect 470 545 476 547
rect 470 543 472 545
rect 474 543 476 545
rect 470 541 476 543
rect 480 546 492 548
rect 497 552 499 561
rect 497 550 503 552
rect 497 548 499 550
rect 501 548 503 550
rect 497 546 503 548
rect 440 530 449 532
rect 443 528 445 530
rect 447 528 449 530
rect 443 526 449 528
rect 473 531 475 541
rect 480 531 482 546
rect 487 540 493 542
rect 487 538 489 540
rect 491 538 493 540
rect 487 536 493 538
rect 490 531 492 536
rect 497 531 499 546
rect 507 543 509 561
rect 539 561 541 566
rect 549 561 551 566
rect 572 572 574 577
rect 579 572 581 577
rect 589 569 591 577
rect 599 569 601 573
rect 612 569 614 577
rect 612 567 617 569
rect 615 564 617 567
rect 529 552 531 555
rect 539 552 541 555
rect 529 550 535 552
rect 529 548 531 550
rect 533 548 535 550
rect 529 546 535 548
rect 539 550 545 552
rect 539 548 541 550
rect 543 548 545 550
rect 539 546 545 548
rect 529 543 531 546
rect 507 532 509 535
rect 507 530 516 532
rect 510 528 512 530
rect 514 528 516 530
rect 510 526 516 528
rect 542 536 544 546
rect 549 545 551 555
rect 572 551 574 560
rect 579 557 581 560
rect 579 555 583 557
rect 589 556 591 560
rect 599 557 601 560
rect 581 552 583 555
rect 599 555 608 557
rect 599 553 604 555
rect 606 553 608 555
rect 571 549 577 551
rect 571 547 573 549
rect 575 547 577 549
rect 571 545 577 547
rect 581 550 587 552
rect 581 548 583 550
rect 585 548 587 550
rect 581 546 587 548
rect 599 551 608 553
rect 599 547 601 551
rect 615 547 617 555
rect 549 543 555 545
rect 549 541 551 543
rect 553 541 555 543
rect 571 542 573 545
rect 581 542 583 546
rect 591 545 601 547
rect 607 545 620 547
rect 591 542 593 545
rect 607 542 609 545
rect 618 544 620 545
rect 618 542 624 544
rect 549 539 555 541
rect 549 536 551 539
rect 529 520 531 525
rect 339 511 341 515
rect 346 511 348 515
rect 356 511 358 515
rect 363 511 365 515
rect 373 511 375 515
rect 396 511 398 515
rect 406 511 408 515
rect 413 511 415 515
rect 423 511 425 515
rect 430 511 432 515
rect 463 511 465 515
rect 473 511 475 515
rect 480 511 482 515
rect 490 511 492 515
rect 497 511 499 515
rect 581 520 583 524
rect 591 520 593 524
rect 542 511 544 515
rect 549 511 551 515
rect 571 511 573 515
rect 618 540 620 542
rect 622 540 624 542
rect 618 538 624 540
rect 607 511 609 515
rect 26 503 28 507
rect 33 503 35 507
rect 13 493 15 498
rect 110 503 112 507
rect 62 494 64 498
rect 72 496 74 501
rect 82 496 84 501
rect 13 472 15 475
rect 26 472 28 482
rect 33 479 35 482
rect 33 477 39 479
rect 33 475 35 477
rect 37 475 39 477
rect 33 473 39 475
rect 13 470 19 472
rect 13 468 15 470
rect 17 468 19 470
rect 13 466 19 468
rect 23 470 29 472
rect 23 468 25 470
rect 27 468 29 470
rect 23 466 29 468
rect 13 463 15 466
rect 23 463 25 466
rect 33 463 35 473
rect 62 472 64 476
rect 72 472 74 483
rect 82 480 84 483
rect 82 478 88 480
rect 82 476 84 478
rect 86 476 88 478
rect 82 474 88 476
rect 95 478 101 480
rect 95 476 97 478
rect 99 476 101 478
rect 146 503 148 507
rect 126 494 128 498
rect 136 494 138 498
rect 224 503 226 507
rect 176 494 178 498
rect 186 496 188 501
rect 196 496 198 501
rect 95 474 101 476
rect 62 470 68 472
rect 62 468 64 470
rect 66 468 68 470
rect 62 466 68 468
rect 72 470 78 472
rect 72 468 74 470
rect 76 468 78 470
rect 72 466 78 468
rect 62 461 64 466
rect 75 461 77 466
rect 82 461 84 474
rect 99 473 101 474
rect 110 473 112 476
rect 126 473 128 476
rect 99 471 112 473
rect 118 471 128 473
rect 136 472 138 476
rect 146 473 148 476
rect 102 463 104 471
rect 118 467 120 471
rect 111 465 120 467
rect 132 470 138 472
rect 132 468 134 470
rect 136 468 138 470
rect 132 466 138 468
rect 142 471 148 473
rect 142 469 144 471
rect 146 469 148 471
rect 142 467 148 469
rect 176 472 178 476
rect 186 472 188 483
rect 196 480 198 483
rect 196 478 202 480
rect 196 476 198 478
rect 200 476 202 478
rect 196 474 202 476
rect 209 478 215 480
rect 209 476 211 478
rect 213 476 215 478
rect 260 503 262 507
rect 240 494 242 498
rect 250 494 252 498
rect 339 503 341 507
rect 346 503 348 507
rect 356 503 358 507
rect 363 503 365 507
rect 373 503 375 507
rect 396 503 398 507
rect 406 503 408 507
rect 413 503 415 507
rect 423 503 425 507
rect 430 503 432 507
rect 463 503 465 507
rect 473 503 475 507
rect 480 503 482 507
rect 490 503 492 507
rect 497 503 499 507
rect 287 496 289 501
rect 297 496 299 501
rect 307 494 309 498
rect 287 480 289 483
rect 283 478 289 480
rect 283 476 285 478
rect 287 476 289 478
rect 209 474 215 476
rect 176 470 182 472
rect 176 468 178 470
rect 180 468 182 470
rect 111 463 113 465
rect 115 463 120 465
rect 13 449 15 454
rect 23 452 25 457
rect 33 452 35 457
rect 62 448 64 452
rect 111 461 120 463
rect 136 463 138 466
rect 118 458 120 461
rect 128 458 130 462
rect 136 461 140 463
rect 138 458 140 461
rect 145 458 147 467
rect 176 466 182 468
rect 186 470 192 472
rect 186 468 188 470
rect 190 468 192 470
rect 186 466 192 468
rect 176 461 178 466
rect 189 461 191 466
rect 196 461 198 474
rect 213 473 215 474
rect 224 473 226 476
rect 240 473 242 476
rect 213 471 226 473
rect 232 471 242 473
rect 250 472 252 476
rect 260 473 262 476
rect 283 474 289 476
rect 216 463 218 471
rect 232 467 234 471
rect 225 465 234 467
rect 246 470 252 472
rect 246 468 248 470
rect 250 468 252 470
rect 246 466 252 468
rect 256 471 262 473
rect 256 469 258 471
rect 260 469 262 471
rect 256 467 262 469
rect 225 463 227 465
rect 229 463 234 465
rect 102 451 104 454
rect 75 445 77 450
rect 82 445 84 450
rect 102 449 107 451
rect 105 441 107 449
rect 118 445 120 449
rect 128 441 130 449
rect 176 448 178 452
rect 225 461 234 463
rect 250 463 252 466
rect 232 458 234 461
rect 242 458 244 462
rect 250 461 254 463
rect 252 458 254 461
rect 259 458 261 467
rect 287 461 289 474
rect 297 472 299 483
rect 322 490 328 492
rect 322 488 324 490
rect 326 488 328 490
rect 322 486 331 488
rect 329 483 331 486
rect 307 472 309 476
rect 293 470 299 472
rect 293 468 295 470
rect 297 468 299 470
rect 293 466 299 468
rect 303 470 309 472
rect 303 468 305 470
rect 307 468 309 470
rect 303 466 309 468
rect 294 461 296 466
rect 307 461 309 466
rect 216 451 218 454
rect 138 441 140 446
rect 145 441 147 446
rect 105 439 130 441
rect 189 445 191 450
rect 196 445 198 450
rect 216 449 221 451
rect 219 441 221 449
rect 232 445 234 449
rect 242 441 244 449
rect 329 457 331 475
rect 339 472 341 487
rect 346 482 348 487
rect 345 480 351 482
rect 345 478 347 480
rect 349 478 351 480
rect 345 476 351 478
rect 356 472 358 487
rect 363 477 365 487
rect 443 490 449 492
rect 443 488 445 490
rect 447 488 449 490
rect 335 470 341 472
rect 335 468 337 470
rect 339 468 341 470
rect 335 466 341 468
rect 339 457 341 466
rect 346 470 358 472
rect 362 475 368 477
rect 362 473 364 475
rect 366 473 368 475
rect 362 471 368 473
rect 346 457 348 470
rect 352 464 358 466
rect 352 462 354 464
rect 356 462 358 464
rect 352 460 358 462
rect 356 457 358 460
rect 363 457 365 471
rect 373 467 375 485
rect 396 467 398 485
rect 406 477 408 487
rect 403 475 409 477
rect 403 473 405 475
rect 407 473 409 475
rect 403 471 409 473
rect 413 472 415 487
rect 423 482 425 487
rect 420 480 426 482
rect 420 478 422 480
rect 424 478 426 480
rect 420 476 426 478
rect 430 472 432 487
rect 440 486 449 488
rect 440 483 442 486
rect 542 503 544 507
rect 549 503 551 507
rect 571 503 573 507
rect 529 493 531 498
rect 510 490 516 492
rect 510 488 512 490
rect 514 488 516 490
rect 370 465 376 467
rect 370 463 372 465
rect 374 463 376 465
rect 370 461 376 463
rect 395 465 401 467
rect 395 463 397 465
rect 399 463 401 465
rect 395 461 401 463
rect 373 458 375 461
rect 396 458 398 461
rect 252 441 254 446
rect 259 441 261 446
rect 287 445 289 450
rect 294 445 296 450
rect 219 439 244 441
rect 307 448 309 452
rect 329 441 331 451
rect 406 457 408 471
rect 413 470 425 472
rect 413 464 419 466
rect 413 462 415 464
rect 417 462 419 464
rect 413 460 419 462
rect 413 457 415 460
rect 423 457 425 470
rect 430 470 436 472
rect 430 468 432 470
rect 434 468 436 470
rect 430 466 436 468
rect 430 457 432 466
rect 440 457 442 475
rect 463 467 465 485
rect 473 477 475 487
rect 470 475 476 477
rect 470 473 472 475
rect 474 473 476 475
rect 470 471 476 473
rect 480 472 482 487
rect 490 482 492 487
rect 487 480 493 482
rect 487 478 489 480
rect 491 478 493 480
rect 487 476 493 478
rect 497 472 499 487
rect 507 486 516 488
rect 507 483 509 486
rect 462 465 468 467
rect 462 463 464 465
rect 466 463 468 465
rect 462 461 468 463
rect 463 458 465 461
rect 339 445 341 449
rect 346 441 348 449
rect 356 444 358 449
rect 363 444 365 449
rect 373 444 375 449
rect 396 444 398 449
rect 406 444 408 449
rect 413 444 415 449
rect 329 439 348 441
rect 423 441 425 449
rect 430 445 432 449
rect 440 441 442 451
rect 473 457 475 471
rect 480 470 492 472
rect 480 464 486 466
rect 480 462 482 464
rect 484 462 486 464
rect 480 460 486 462
rect 480 457 482 460
rect 490 457 492 470
rect 497 470 503 472
rect 497 468 499 470
rect 501 468 503 470
rect 497 466 503 468
rect 497 457 499 466
rect 507 457 509 475
rect 529 472 531 475
rect 542 472 544 482
rect 549 479 551 482
rect 549 477 555 479
rect 549 475 551 477
rect 553 475 555 477
rect 607 503 609 507
rect 581 494 583 498
rect 591 494 593 498
rect 618 478 624 480
rect 618 476 620 478
rect 622 476 624 478
rect 549 473 555 475
rect 571 473 573 476
rect 529 470 535 472
rect 529 468 531 470
rect 533 468 535 470
rect 529 466 535 468
rect 539 470 545 472
rect 539 468 541 470
rect 543 468 545 470
rect 539 466 545 468
rect 529 463 531 466
rect 539 463 541 466
rect 549 463 551 473
rect 571 471 577 473
rect 571 469 573 471
rect 575 469 577 471
rect 571 467 577 469
rect 581 472 583 476
rect 591 473 593 476
rect 607 473 609 476
rect 618 474 624 476
rect 618 473 620 474
rect 581 470 587 472
rect 591 471 601 473
rect 607 471 620 473
rect 581 468 583 470
rect 585 468 587 470
rect 572 458 574 467
rect 581 466 587 468
rect 599 467 601 471
rect 581 463 583 466
rect 579 461 583 463
rect 599 465 608 467
rect 599 463 604 465
rect 606 463 608 465
rect 615 463 617 471
rect 579 458 581 461
rect 589 458 591 462
rect 599 461 608 463
rect 599 458 601 461
rect 463 444 465 449
rect 473 444 475 449
rect 480 444 482 449
rect 423 439 442 441
rect 490 441 492 449
rect 497 445 499 449
rect 507 441 509 451
rect 529 449 531 454
rect 539 452 541 457
rect 549 452 551 457
rect 490 439 509 441
rect 615 451 617 454
rect 612 449 617 451
rect 572 441 574 446
rect 579 441 581 446
rect 589 441 591 449
rect 599 445 601 449
rect 612 441 614 449
rect 589 439 614 441
rect 13 420 15 425
rect 23 417 25 422
rect 33 417 35 422
rect 62 422 64 426
rect 75 424 77 429
rect 82 424 84 429
rect 105 433 130 435
rect 105 425 107 433
rect 118 425 120 429
rect 128 425 130 433
rect 138 428 140 433
rect 145 428 147 433
rect 102 423 107 425
rect 102 420 104 423
rect 13 408 15 411
rect 23 408 25 411
rect 13 406 19 408
rect 13 404 15 406
rect 17 404 19 406
rect 13 402 19 404
rect 23 406 29 408
rect 23 404 25 406
rect 27 404 29 406
rect 23 402 29 404
rect 13 399 15 402
rect 26 392 28 402
rect 33 401 35 411
rect 62 408 64 413
rect 75 408 77 413
rect 62 406 68 408
rect 62 404 64 406
rect 66 404 68 406
rect 62 402 68 404
rect 72 406 78 408
rect 72 404 74 406
rect 76 404 78 406
rect 72 402 78 404
rect 33 399 39 401
rect 33 397 35 399
rect 37 397 39 399
rect 62 398 64 402
rect 33 395 39 397
rect 33 392 35 395
rect 13 376 15 381
rect 72 391 74 402
rect 82 400 84 413
rect 176 422 178 426
rect 189 424 191 429
rect 196 424 198 429
rect 219 433 244 435
rect 219 425 221 433
rect 232 425 234 429
rect 242 425 244 433
rect 252 428 254 433
rect 259 428 261 433
rect 118 413 120 416
rect 111 411 120 413
rect 128 412 130 416
rect 138 413 140 416
rect 102 403 104 411
rect 111 409 113 411
rect 115 409 120 411
rect 111 407 120 409
rect 136 411 140 413
rect 136 408 138 411
rect 118 403 120 407
rect 132 406 138 408
rect 145 407 147 416
rect 216 423 221 425
rect 216 420 218 423
rect 176 408 178 413
rect 189 408 191 413
rect 132 404 134 406
rect 136 404 138 406
rect 99 401 112 403
rect 118 401 128 403
rect 132 402 138 404
rect 99 400 101 401
rect 82 398 88 400
rect 82 396 84 398
rect 86 396 88 398
rect 82 394 88 396
rect 95 398 101 400
rect 110 398 112 401
rect 126 398 128 401
rect 136 398 138 402
rect 142 405 148 407
rect 142 403 144 405
rect 146 403 148 405
rect 142 401 148 403
rect 146 398 148 401
rect 176 406 182 408
rect 176 404 178 406
rect 180 404 182 406
rect 176 402 182 404
rect 186 406 192 408
rect 186 404 188 406
rect 190 404 192 406
rect 186 402 192 404
rect 176 398 178 402
rect 95 396 97 398
rect 99 396 101 398
rect 95 394 101 396
rect 82 391 84 394
rect 62 376 64 380
rect 72 373 74 378
rect 82 373 84 378
rect 26 367 28 371
rect 33 367 35 371
rect 126 376 128 380
rect 136 376 138 380
rect 110 367 112 371
rect 186 391 188 402
rect 196 400 198 413
rect 287 424 289 429
rect 294 424 296 429
rect 329 433 348 435
rect 232 413 234 416
rect 225 411 234 413
rect 242 412 244 416
rect 252 413 254 416
rect 216 403 218 411
rect 225 409 227 411
rect 229 409 234 411
rect 225 407 234 409
rect 250 411 254 413
rect 250 408 252 411
rect 232 403 234 407
rect 246 406 252 408
rect 259 407 261 416
rect 307 422 309 426
rect 329 423 331 433
rect 339 425 341 429
rect 346 425 348 433
rect 423 433 442 435
rect 356 425 358 430
rect 363 425 365 430
rect 373 425 375 430
rect 396 425 398 430
rect 406 425 408 430
rect 413 425 415 430
rect 423 425 425 433
rect 430 425 432 429
rect 246 404 248 406
rect 250 404 252 406
rect 213 401 226 403
rect 232 401 242 403
rect 246 402 252 404
rect 213 400 215 401
rect 196 398 202 400
rect 196 396 198 398
rect 200 396 202 398
rect 196 394 202 396
rect 209 398 215 400
rect 224 398 226 401
rect 240 398 242 401
rect 250 398 252 402
rect 256 405 262 407
rect 256 403 258 405
rect 260 403 262 405
rect 256 401 262 403
rect 260 398 262 401
rect 287 400 289 413
rect 294 408 296 413
rect 307 408 309 413
rect 293 406 299 408
rect 293 404 295 406
rect 297 404 299 406
rect 293 402 299 404
rect 303 406 309 408
rect 303 404 305 406
rect 307 404 309 406
rect 303 402 309 404
rect 283 398 289 400
rect 209 396 211 398
rect 213 396 215 398
rect 209 394 215 396
rect 196 391 198 394
rect 176 376 178 380
rect 186 373 188 378
rect 196 373 198 378
rect 146 367 148 371
rect 240 376 242 380
rect 250 376 252 380
rect 224 367 226 371
rect 283 396 285 398
rect 287 396 289 398
rect 283 394 289 396
rect 287 391 289 394
rect 297 391 299 402
rect 307 398 309 402
rect 329 399 331 417
rect 339 408 341 417
rect 335 406 341 408
rect 335 404 337 406
rect 339 404 341 406
rect 335 402 341 404
rect 346 404 348 417
rect 356 414 358 417
rect 352 412 358 414
rect 352 410 354 412
rect 356 410 358 412
rect 352 408 358 410
rect 346 402 358 404
rect 363 403 365 417
rect 440 423 442 433
rect 490 433 509 435
rect 463 425 465 430
rect 473 425 475 430
rect 480 425 482 430
rect 490 425 492 433
rect 497 425 499 429
rect 373 413 375 416
rect 396 413 398 416
rect 370 411 376 413
rect 370 409 372 411
rect 374 409 376 411
rect 370 407 376 409
rect 395 411 401 413
rect 395 409 397 411
rect 399 409 401 411
rect 395 407 401 409
rect 329 388 331 391
rect 322 386 331 388
rect 339 387 341 402
rect 345 396 351 398
rect 345 394 347 396
rect 349 394 351 396
rect 345 392 351 394
rect 346 387 348 392
rect 356 387 358 402
rect 362 401 368 403
rect 362 399 364 401
rect 366 399 368 401
rect 362 397 368 399
rect 363 387 365 397
rect 373 389 375 407
rect 396 389 398 407
rect 406 403 408 417
rect 413 414 415 417
rect 413 412 419 414
rect 413 410 415 412
rect 417 410 419 412
rect 413 408 419 410
rect 423 404 425 417
rect 403 401 409 403
rect 403 399 405 401
rect 407 399 409 401
rect 403 397 409 399
rect 413 402 425 404
rect 430 408 432 417
rect 430 406 436 408
rect 430 404 432 406
rect 434 404 436 406
rect 430 402 436 404
rect 322 384 324 386
rect 326 384 328 386
rect 322 382 328 384
rect 287 373 289 378
rect 297 373 299 378
rect 307 376 309 380
rect 260 367 262 371
rect 406 387 408 397
rect 413 387 415 402
rect 420 396 426 398
rect 420 394 422 396
rect 424 394 426 396
rect 420 392 426 394
rect 423 387 425 392
rect 430 387 432 402
rect 440 399 442 417
rect 507 423 509 433
rect 589 433 614 435
rect 529 420 531 425
rect 463 413 465 416
rect 462 411 468 413
rect 462 409 464 411
rect 466 409 468 411
rect 462 407 468 409
rect 440 388 442 391
rect 463 389 465 407
rect 473 403 475 417
rect 480 414 482 417
rect 480 412 486 414
rect 480 410 482 412
rect 484 410 486 412
rect 480 408 486 410
rect 490 404 492 417
rect 470 401 476 403
rect 470 399 472 401
rect 474 399 476 401
rect 470 397 476 399
rect 480 402 492 404
rect 497 408 499 417
rect 497 406 503 408
rect 497 404 499 406
rect 501 404 503 406
rect 497 402 503 404
rect 440 386 449 388
rect 443 384 445 386
rect 447 384 449 386
rect 443 382 449 384
rect 473 387 475 397
rect 480 387 482 402
rect 487 396 493 398
rect 487 394 489 396
rect 491 394 493 396
rect 487 392 493 394
rect 490 387 492 392
rect 497 387 499 402
rect 507 399 509 417
rect 539 417 541 422
rect 549 417 551 422
rect 572 428 574 433
rect 579 428 581 433
rect 589 425 591 433
rect 599 425 601 429
rect 612 425 614 433
rect 612 423 617 425
rect 615 420 617 423
rect 529 408 531 411
rect 539 408 541 411
rect 529 406 535 408
rect 529 404 531 406
rect 533 404 535 406
rect 529 402 535 404
rect 539 406 545 408
rect 539 404 541 406
rect 543 404 545 406
rect 539 402 545 404
rect 529 399 531 402
rect 507 388 509 391
rect 507 386 516 388
rect 510 384 512 386
rect 514 384 516 386
rect 510 382 516 384
rect 542 392 544 402
rect 549 401 551 411
rect 572 407 574 416
rect 579 413 581 416
rect 579 411 583 413
rect 589 412 591 416
rect 599 413 601 416
rect 581 408 583 411
rect 599 411 608 413
rect 599 409 604 411
rect 606 409 608 411
rect 571 405 577 407
rect 571 403 573 405
rect 575 403 577 405
rect 571 401 577 403
rect 581 406 587 408
rect 581 404 583 406
rect 585 404 587 406
rect 581 402 587 404
rect 599 407 608 409
rect 599 403 601 407
rect 615 403 617 411
rect 549 399 555 401
rect 549 397 551 399
rect 553 397 555 399
rect 571 398 573 401
rect 581 398 583 402
rect 591 401 601 403
rect 607 401 620 403
rect 591 398 593 401
rect 607 398 609 401
rect 618 400 620 401
rect 618 398 624 400
rect 549 395 555 397
rect 549 392 551 395
rect 529 376 531 381
rect 339 367 341 371
rect 346 367 348 371
rect 356 367 358 371
rect 363 367 365 371
rect 373 367 375 371
rect 396 367 398 371
rect 406 367 408 371
rect 413 367 415 371
rect 423 367 425 371
rect 430 367 432 371
rect 463 367 465 371
rect 473 367 475 371
rect 480 367 482 371
rect 490 367 492 371
rect 497 367 499 371
rect 581 376 583 380
rect 591 376 593 380
rect 542 367 544 371
rect 549 367 551 371
rect 571 367 573 371
rect 618 396 620 398
rect 622 396 624 398
rect 618 394 624 396
rect 607 367 609 371
rect 26 359 28 363
rect 33 359 35 363
rect 13 349 15 354
rect 110 359 112 363
rect 62 350 64 354
rect 72 352 74 357
rect 82 352 84 357
rect 13 328 15 331
rect 26 328 28 338
rect 33 335 35 338
rect 33 333 39 335
rect 33 331 35 333
rect 37 331 39 333
rect 33 329 39 331
rect 13 326 19 328
rect 13 324 15 326
rect 17 324 19 326
rect 13 322 19 324
rect 23 326 29 328
rect 23 324 25 326
rect 27 324 29 326
rect 23 322 29 324
rect 13 319 15 322
rect 23 319 25 322
rect 33 319 35 329
rect 62 328 64 332
rect 72 328 74 339
rect 82 336 84 339
rect 82 334 88 336
rect 82 332 84 334
rect 86 332 88 334
rect 82 330 88 332
rect 95 334 101 336
rect 95 332 97 334
rect 99 332 101 334
rect 146 359 148 363
rect 126 350 128 354
rect 136 350 138 354
rect 224 359 226 363
rect 176 350 178 354
rect 186 352 188 357
rect 196 352 198 357
rect 95 330 101 332
rect 62 326 68 328
rect 62 324 64 326
rect 66 324 68 326
rect 62 322 68 324
rect 72 326 78 328
rect 72 324 74 326
rect 76 324 78 326
rect 72 322 78 324
rect 62 317 64 322
rect 75 317 77 322
rect 82 317 84 330
rect 99 329 101 330
rect 110 329 112 332
rect 126 329 128 332
rect 99 327 112 329
rect 118 327 128 329
rect 136 328 138 332
rect 146 329 148 332
rect 102 319 104 327
rect 118 323 120 327
rect 111 321 120 323
rect 132 326 138 328
rect 132 324 134 326
rect 136 324 138 326
rect 132 322 138 324
rect 142 327 148 329
rect 142 325 144 327
rect 146 325 148 327
rect 142 323 148 325
rect 176 328 178 332
rect 186 328 188 339
rect 196 336 198 339
rect 196 334 202 336
rect 196 332 198 334
rect 200 332 202 334
rect 196 330 202 332
rect 209 334 215 336
rect 209 332 211 334
rect 213 332 215 334
rect 260 359 262 363
rect 240 350 242 354
rect 250 350 252 354
rect 339 359 341 363
rect 346 359 348 363
rect 356 359 358 363
rect 363 359 365 363
rect 373 359 375 363
rect 396 359 398 363
rect 406 359 408 363
rect 413 359 415 363
rect 423 359 425 363
rect 430 359 432 363
rect 463 359 465 363
rect 473 359 475 363
rect 480 359 482 363
rect 490 359 492 363
rect 497 359 499 363
rect 287 352 289 357
rect 297 352 299 357
rect 307 350 309 354
rect 287 336 289 339
rect 283 334 289 336
rect 283 332 285 334
rect 287 332 289 334
rect 209 330 215 332
rect 176 326 182 328
rect 176 324 178 326
rect 180 324 182 326
rect 111 319 113 321
rect 115 319 120 321
rect 13 305 15 310
rect 23 308 25 313
rect 33 308 35 313
rect 62 304 64 308
rect 111 317 120 319
rect 136 319 138 322
rect 118 314 120 317
rect 128 314 130 318
rect 136 317 140 319
rect 138 314 140 317
rect 145 314 147 323
rect 176 322 182 324
rect 186 326 192 328
rect 186 324 188 326
rect 190 324 192 326
rect 186 322 192 324
rect 176 317 178 322
rect 189 317 191 322
rect 196 317 198 330
rect 213 329 215 330
rect 224 329 226 332
rect 240 329 242 332
rect 213 327 226 329
rect 232 327 242 329
rect 250 328 252 332
rect 260 329 262 332
rect 283 330 289 332
rect 216 319 218 327
rect 232 323 234 327
rect 225 321 234 323
rect 246 326 252 328
rect 246 324 248 326
rect 250 324 252 326
rect 246 322 252 324
rect 256 327 262 329
rect 256 325 258 327
rect 260 325 262 327
rect 256 323 262 325
rect 225 319 227 321
rect 229 319 234 321
rect 102 307 104 310
rect 75 301 77 306
rect 82 301 84 306
rect 102 305 107 307
rect 105 297 107 305
rect 118 301 120 305
rect 128 297 130 305
rect 176 304 178 308
rect 225 317 234 319
rect 250 319 252 322
rect 232 314 234 317
rect 242 314 244 318
rect 250 317 254 319
rect 252 314 254 317
rect 259 314 261 323
rect 287 317 289 330
rect 297 328 299 339
rect 322 346 328 348
rect 322 344 324 346
rect 326 344 328 346
rect 322 342 331 344
rect 329 339 331 342
rect 307 328 309 332
rect 293 326 299 328
rect 293 324 295 326
rect 297 324 299 326
rect 293 322 299 324
rect 303 326 309 328
rect 303 324 305 326
rect 307 324 309 326
rect 303 322 309 324
rect 294 317 296 322
rect 307 317 309 322
rect 216 307 218 310
rect 138 297 140 302
rect 145 297 147 302
rect 105 295 130 297
rect 189 301 191 306
rect 196 301 198 306
rect 216 305 221 307
rect 219 297 221 305
rect 232 301 234 305
rect 242 297 244 305
rect 329 313 331 331
rect 339 328 341 343
rect 346 338 348 343
rect 345 336 351 338
rect 345 334 347 336
rect 349 334 351 336
rect 345 332 351 334
rect 356 328 358 343
rect 363 333 365 343
rect 443 346 449 348
rect 443 344 445 346
rect 447 344 449 346
rect 335 326 341 328
rect 335 324 337 326
rect 339 324 341 326
rect 335 322 341 324
rect 339 313 341 322
rect 346 326 358 328
rect 362 331 368 333
rect 362 329 364 331
rect 366 329 368 331
rect 362 327 368 329
rect 346 313 348 326
rect 352 320 358 322
rect 352 318 354 320
rect 356 318 358 320
rect 352 316 358 318
rect 356 313 358 316
rect 363 313 365 327
rect 373 323 375 341
rect 396 323 398 341
rect 406 333 408 343
rect 403 331 409 333
rect 403 329 405 331
rect 407 329 409 331
rect 403 327 409 329
rect 413 328 415 343
rect 423 338 425 343
rect 420 336 426 338
rect 420 334 422 336
rect 424 334 426 336
rect 420 332 426 334
rect 430 328 432 343
rect 440 342 449 344
rect 440 339 442 342
rect 542 359 544 363
rect 549 359 551 363
rect 571 359 573 363
rect 529 349 531 354
rect 510 346 516 348
rect 510 344 512 346
rect 514 344 516 346
rect 370 321 376 323
rect 370 319 372 321
rect 374 319 376 321
rect 370 317 376 319
rect 395 321 401 323
rect 395 319 397 321
rect 399 319 401 321
rect 395 317 401 319
rect 373 314 375 317
rect 396 314 398 317
rect 252 297 254 302
rect 259 297 261 302
rect 287 301 289 306
rect 294 301 296 306
rect 219 295 244 297
rect 307 304 309 308
rect 329 297 331 307
rect 406 313 408 327
rect 413 326 425 328
rect 413 320 419 322
rect 413 318 415 320
rect 417 318 419 320
rect 413 316 419 318
rect 413 313 415 316
rect 423 313 425 326
rect 430 326 436 328
rect 430 324 432 326
rect 434 324 436 326
rect 430 322 436 324
rect 430 313 432 322
rect 440 313 442 331
rect 463 323 465 341
rect 473 333 475 343
rect 470 331 476 333
rect 470 329 472 331
rect 474 329 476 331
rect 470 327 476 329
rect 480 328 482 343
rect 490 338 492 343
rect 487 336 493 338
rect 487 334 489 336
rect 491 334 493 336
rect 487 332 493 334
rect 497 328 499 343
rect 507 342 516 344
rect 507 339 509 342
rect 462 321 468 323
rect 462 319 464 321
rect 466 319 468 321
rect 462 317 468 319
rect 463 314 465 317
rect 339 301 341 305
rect 346 297 348 305
rect 356 300 358 305
rect 363 300 365 305
rect 373 300 375 305
rect 396 300 398 305
rect 406 300 408 305
rect 413 300 415 305
rect 329 295 348 297
rect 423 297 425 305
rect 430 301 432 305
rect 440 297 442 307
rect 473 313 475 327
rect 480 326 492 328
rect 480 320 486 322
rect 480 318 482 320
rect 484 318 486 320
rect 480 316 486 318
rect 480 313 482 316
rect 490 313 492 326
rect 497 326 503 328
rect 497 324 499 326
rect 501 324 503 326
rect 497 322 503 324
rect 497 313 499 322
rect 507 313 509 331
rect 529 328 531 331
rect 542 328 544 338
rect 549 335 551 338
rect 549 333 555 335
rect 549 331 551 333
rect 553 331 555 333
rect 607 359 609 363
rect 581 350 583 354
rect 591 350 593 354
rect 618 334 624 336
rect 618 332 620 334
rect 622 332 624 334
rect 549 329 555 331
rect 571 329 573 332
rect 529 326 535 328
rect 529 324 531 326
rect 533 324 535 326
rect 529 322 535 324
rect 539 326 545 328
rect 539 324 541 326
rect 543 324 545 326
rect 539 322 545 324
rect 529 319 531 322
rect 539 319 541 322
rect 549 319 551 329
rect 571 327 577 329
rect 571 325 573 327
rect 575 325 577 327
rect 571 323 577 325
rect 581 328 583 332
rect 591 329 593 332
rect 607 329 609 332
rect 618 330 624 332
rect 618 329 620 330
rect 581 326 587 328
rect 591 327 601 329
rect 607 327 620 329
rect 581 324 583 326
rect 585 324 587 326
rect 572 314 574 323
rect 581 322 587 324
rect 599 323 601 327
rect 581 319 583 322
rect 579 317 583 319
rect 599 321 608 323
rect 599 319 604 321
rect 606 319 608 321
rect 615 319 617 327
rect 579 314 581 317
rect 589 314 591 318
rect 599 317 608 319
rect 599 314 601 317
rect 463 300 465 305
rect 473 300 475 305
rect 480 300 482 305
rect 423 295 442 297
rect 490 297 492 305
rect 497 301 499 305
rect 507 297 509 307
rect 529 305 531 310
rect 539 308 541 313
rect 549 308 551 313
rect 490 295 509 297
rect 615 307 617 310
rect 612 305 617 307
rect 572 297 574 302
rect 579 297 581 302
rect 589 297 591 305
rect 599 301 601 305
rect 612 297 614 305
rect 589 295 614 297
rect 13 276 15 281
rect 23 273 25 278
rect 33 273 35 278
rect 62 278 64 282
rect 75 280 77 285
rect 82 280 84 285
rect 105 289 130 291
rect 105 281 107 289
rect 118 281 120 285
rect 128 281 130 289
rect 138 284 140 289
rect 145 284 147 289
rect 102 279 107 281
rect 102 276 104 279
rect 13 264 15 267
rect 23 264 25 267
rect 13 262 19 264
rect 13 260 15 262
rect 17 260 19 262
rect 13 258 19 260
rect 23 262 29 264
rect 23 260 25 262
rect 27 260 29 262
rect 23 258 29 260
rect 13 255 15 258
rect 26 248 28 258
rect 33 257 35 267
rect 62 264 64 269
rect 75 264 77 269
rect 62 262 68 264
rect 62 260 64 262
rect 66 260 68 262
rect 62 258 68 260
rect 72 262 78 264
rect 72 260 74 262
rect 76 260 78 262
rect 72 258 78 260
rect 33 255 39 257
rect 33 253 35 255
rect 37 253 39 255
rect 62 254 64 258
rect 33 251 39 253
rect 33 248 35 251
rect 13 232 15 237
rect 72 247 74 258
rect 82 256 84 269
rect 176 278 178 282
rect 189 280 191 285
rect 196 280 198 285
rect 219 289 244 291
rect 219 281 221 289
rect 232 281 234 285
rect 242 281 244 289
rect 252 284 254 289
rect 259 284 261 289
rect 118 269 120 272
rect 111 267 120 269
rect 128 268 130 272
rect 138 269 140 272
rect 102 259 104 267
rect 111 265 113 267
rect 115 265 120 267
rect 111 263 120 265
rect 136 267 140 269
rect 136 264 138 267
rect 118 259 120 263
rect 132 262 138 264
rect 145 263 147 272
rect 216 279 221 281
rect 216 276 218 279
rect 176 264 178 269
rect 189 264 191 269
rect 132 260 134 262
rect 136 260 138 262
rect 99 257 112 259
rect 118 257 128 259
rect 132 258 138 260
rect 99 256 101 257
rect 82 254 88 256
rect 82 252 84 254
rect 86 252 88 254
rect 82 250 88 252
rect 95 254 101 256
rect 110 254 112 257
rect 126 254 128 257
rect 136 254 138 258
rect 142 261 148 263
rect 142 259 144 261
rect 146 259 148 261
rect 142 257 148 259
rect 146 254 148 257
rect 176 262 182 264
rect 176 260 178 262
rect 180 260 182 262
rect 176 258 182 260
rect 186 262 192 264
rect 186 260 188 262
rect 190 260 192 262
rect 186 258 192 260
rect 176 254 178 258
rect 95 252 97 254
rect 99 252 101 254
rect 95 250 101 252
rect 82 247 84 250
rect 62 232 64 236
rect 72 229 74 234
rect 82 229 84 234
rect 26 223 28 227
rect 33 223 35 227
rect 126 232 128 236
rect 136 232 138 236
rect 110 223 112 227
rect 186 247 188 258
rect 196 256 198 269
rect 287 280 289 285
rect 294 280 296 285
rect 329 289 348 291
rect 232 269 234 272
rect 225 267 234 269
rect 242 268 244 272
rect 252 269 254 272
rect 216 259 218 267
rect 225 265 227 267
rect 229 265 234 267
rect 225 263 234 265
rect 250 267 254 269
rect 250 264 252 267
rect 232 259 234 263
rect 246 262 252 264
rect 259 263 261 272
rect 307 278 309 282
rect 329 279 331 289
rect 339 281 341 285
rect 346 281 348 289
rect 423 289 442 291
rect 356 281 358 286
rect 363 281 365 286
rect 373 281 375 286
rect 396 281 398 286
rect 406 281 408 286
rect 413 281 415 286
rect 423 281 425 289
rect 430 281 432 285
rect 246 260 248 262
rect 250 260 252 262
rect 213 257 226 259
rect 232 257 242 259
rect 246 258 252 260
rect 213 256 215 257
rect 196 254 202 256
rect 196 252 198 254
rect 200 252 202 254
rect 196 250 202 252
rect 209 254 215 256
rect 224 254 226 257
rect 240 254 242 257
rect 250 254 252 258
rect 256 261 262 263
rect 256 259 258 261
rect 260 259 262 261
rect 256 257 262 259
rect 260 254 262 257
rect 287 256 289 269
rect 294 264 296 269
rect 307 264 309 269
rect 293 262 299 264
rect 293 260 295 262
rect 297 260 299 262
rect 293 258 299 260
rect 303 262 309 264
rect 303 260 305 262
rect 307 260 309 262
rect 303 258 309 260
rect 283 254 289 256
rect 209 252 211 254
rect 213 252 215 254
rect 209 250 215 252
rect 196 247 198 250
rect 176 232 178 236
rect 186 229 188 234
rect 196 229 198 234
rect 146 223 148 227
rect 240 232 242 236
rect 250 232 252 236
rect 224 223 226 227
rect 283 252 285 254
rect 287 252 289 254
rect 283 250 289 252
rect 287 247 289 250
rect 297 247 299 258
rect 307 254 309 258
rect 329 255 331 273
rect 339 264 341 273
rect 335 262 341 264
rect 335 260 337 262
rect 339 260 341 262
rect 335 258 341 260
rect 346 260 348 273
rect 356 270 358 273
rect 352 268 358 270
rect 352 266 354 268
rect 356 266 358 268
rect 352 264 358 266
rect 346 258 358 260
rect 363 259 365 273
rect 440 279 442 289
rect 490 289 509 291
rect 463 281 465 286
rect 473 281 475 286
rect 480 281 482 286
rect 490 281 492 289
rect 497 281 499 285
rect 373 269 375 272
rect 396 269 398 272
rect 370 267 376 269
rect 370 265 372 267
rect 374 265 376 267
rect 370 263 376 265
rect 395 267 401 269
rect 395 265 397 267
rect 399 265 401 267
rect 395 263 401 265
rect 329 244 331 247
rect 322 242 331 244
rect 339 243 341 258
rect 345 252 351 254
rect 345 250 347 252
rect 349 250 351 252
rect 345 248 351 250
rect 346 243 348 248
rect 356 243 358 258
rect 362 257 368 259
rect 362 255 364 257
rect 366 255 368 257
rect 362 253 368 255
rect 363 243 365 253
rect 373 245 375 263
rect 396 245 398 263
rect 406 259 408 273
rect 413 270 415 273
rect 413 268 419 270
rect 413 266 415 268
rect 417 266 419 268
rect 413 264 419 266
rect 423 260 425 273
rect 403 257 409 259
rect 403 255 405 257
rect 407 255 409 257
rect 403 253 409 255
rect 413 258 425 260
rect 430 264 432 273
rect 430 262 436 264
rect 430 260 432 262
rect 434 260 436 262
rect 430 258 436 260
rect 322 240 324 242
rect 326 240 328 242
rect 322 238 328 240
rect 287 229 289 234
rect 297 229 299 234
rect 307 232 309 236
rect 260 223 262 227
rect 406 243 408 253
rect 413 243 415 258
rect 420 252 426 254
rect 420 250 422 252
rect 424 250 426 252
rect 420 248 426 250
rect 423 243 425 248
rect 430 243 432 258
rect 440 255 442 273
rect 507 279 509 289
rect 589 289 614 291
rect 529 276 531 281
rect 463 269 465 272
rect 462 267 468 269
rect 462 265 464 267
rect 466 265 468 267
rect 462 263 468 265
rect 440 244 442 247
rect 463 245 465 263
rect 473 259 475 273
rect 480 270 482 273
rect 480 268 486 270
rect 480 266 482 268
rect 484 266 486 268
rect 480 264 486 266
rect 490 260 492 273
rect 470 257 476 259
rect 470 255 472 257
rect 474 255 476 257
rect 470 253 476 255
rect 480 258 492 260
rect 497 264 499 273
rect 497 262 503 264
rect 497 260 499 262
rect 501 260 503 262
rect 497 258 503 260
rect 440 242 449 244
rect 443 240 445 242
rect 447 240 449 242
rect 443 238 449 240
rect 473 243 475 253
rect 480 243 482 258
rect 487 252 493 254
rect 487 250 489 252
rect 491 250 493 252
rect 487 248 493 250
rect 490 243 492 248
rect 497 243 499 258
rect 507 255 509 273
rect 539 273 541 278
rect 549 273 551 278
rect 572 284 574 289
rect 579 284 581 289
rect 589 281 591 289
rect 599 281 601 285
rect 612 281 614 289
rect 612 279 617 281
rect 615 276 617 279
rect 529 264 531 267
rect 539 264 541 267
rect 529 262 535 264
rect 529 260 531 262
rect 533 260 535 262
rect 529 258 535 260
rect 539 262 545 264
rect 539 260 541 262
rect 543 260 545 262
rect 539 258 545 260
rect 529 255 531 258
rect 507 244 509 247
rect 507 242 516 244
rect 510 240 512 242
rect 514 240 516 242
rect 510 238 516 240
rect 542 248 544 258
rect 549 257 551 267
rect 572 263 574 272
rect 579 269 581 272
rect 579 267 583 269
rect 589 268 591 272
rect 599 269 601 272
rect 581 264 583 267
rect 599 267 608 269
rect 599 265 604 267
rect 606 265 608 267
rect 571 261 577 263
rect 571 259 573 261
rect 575 259 577 261
rect 571 257 577 259
rect 581 262 587 264
rect 581 260 583 262
rect 585 260 587 262
rect 581 258 587 260
rect 599 263 608 265
rect 599 259 601 263
rect 615 259 617 267
rect 549 255 555 257
rect 549 253 551 255
rect 553 253 555 255
rect 571 254 573 257
rect 581 254 583 258
rect 591 257 601 259
rect 607 257 620 259
rect 591 254 593 257
rect 607 254 609 257
rect 618 256 620 257
rect 618 254 624 256
rect 549 251 555 253
rect 549 248 551 251
rect 529 232 531 237
rect 339 223 341 227
rect 346 223 348 227
rect 356 223 358 227
rect 363 223 365 227
rect 373 223 375 227
rect 396 223 398 227
rect 406 223 408 227
rect 413 223 415 227
rect 423 223 425 227
rect 430 223 432 227
rect 463 223 465 227
rect 473 223 475 227
rect 480 223 482 227
rect 490 223 492 227
rect 497 223 499 227
rect 581 232 583 236
rect 591 232 593 236
rect 542 223 544 227
rect 549 223 551 227
rect 571 223 573 227
rect 618 252 620 254
rect 622 252 624 254
rect 618 250 624 252
rect 607 223 609 227
rect 26 215 28 219
rect 33 215 35 219
rect 13 205 15 210
rect 110 215 112 219
rect 62 206 64 210
rect 72 208 74 213
rect 82 208 84 213
rect 13 184 15 187
rect 26 184 28 194
rect 33 191 35 194
rect 33 189 39 191
rect 33 187 35 189
rect 37 187 39 189
rect 33 185 39 187
rect 13 182 19 184
rect 13 180 15 182
rect 17 180 19 182
rect 13 178 19 180
rect 23 182 29 184
rect 23 180 25 182
rect 27 180 29 182
rect 23 178 29 180
rect 13 175 15 178
rect 23 175 25 178
rect 33 175 35 185
rect 62 184 64 188
rect 72 184 74 195
rect 82 192 84 195
rect 82 190 88 192
rect 82 188 84 190
rect 86 188 88 190
rect 82 186 88 188
rect 95 190 101 192
rect 95 188 97 190
rect 99 188 101 190
rect 146 215 148 219
rect 126 206 128 210
rect 136 206 138 210
rect 224 215 226 219
rect 176 206 178 210
rect 186 208 188 213
rect 196 208 198 213
rect 95 186 101 188
rect 62 182 68 184
rect 62 180 64 182
rect 66 180 68 182
rect 62 178 68 180
rect 72 182 78 184
rect 72 180 74 182
rect 76 180 78 182
rect 72 178 78 180
rect 62 173 64 178
rect 75 173 77 178
rect 82 173 84 186
rect 99 185 101 186
rect 110 185 112 188
rect 126 185 128 188
rect 99 183 112 185
rect 118 183 128 185
rect 136 184 138 188
rect 146 185 148 188
rect 102 175 104 183
rect 118 179 120 183
rect 111 177 120 179
rect 132 182 138 184
rect 132 180 134 182
rect 136 180 138 182
rect 132 178 138 180
rect 142 183 148 185
rect 142 181 144 183
rect 146 181 148 183
rect 142 179 148 181
rect 176 184 178 188
rect 186 184 188 195
rect 196 192 198 195
rect 196 190 202 192
rect 196 188 198 190
rect 200 188 202 190
rect 196 186 202 188
rect 209 190 215 192
rect 209 188 211 190
rect 213 188 215 190
rect 260 215 262 219
rect 240 206 242 210
rect 250 206 252 210
rect 339 215 341 219
rect 346 215 348 219
rect 356 215 358 219
rect 363 215 365 219
rect 373 215 375 219
rect 396 215 398 219
rect 406 215 408 219
rect 413 215 415 219
rect 423 215 425 219
rect 430 215 432 219
rect 463 215 465 219
rect 473 215 475 219
rect 480 215 482 219
rect 490 215 492 219
rect 497 215 499 219
rect 287 208 289 213
rect 297 208 299 213
rect 307 206 309 210
rect 287 192 289 195
rect 283 190 289 192
rect 283 188 285 190
rect 287 188 289 190
rect 209 186 215 188
rect 176 182 182 184
rect 176 180 178 182
rect 180 180 182 182
rect 111 175 113 177
rect 115 175 120 177
rect 13 161 15 166
rect 23 164 25 169
rect 33 164 35 169
rect 62 160 64 164
rect 111 173 120 175
rect 136 175 138 178
rect 118 170 120 173
rect 128 170 130 174
rect 136 173 140 175
rect 138 170 140 173
rect 145 170 147 179
rect 176 178 182 180
rect 186 182 192 184
rect 186 180 188 182
rect 190 180 192 182
rect 186 178 192 180
rect 176 173 178 178
rect 189 173 191 178
rect 196 173 198 186
rect 213 185 215 186
rect 224 185 226 188
rect 240 185 242 188
rect 213 183 226 185
rect 232 183 242 185
rect 250 184 252 188
rect 260 185 262 188
rect 283 186 289 188
rect 216 175 218 183
rect 232 179 234 183
rect 225 177 234 179
rect 246 182 252 184
rect 246 180 248 182
rect 250 180 252 182
rect 246 178 252 180
rect 256 183 262 185
rect 256 181 258 183
rect 260 181 262 183
rect 256 179 262 181
rect 225 175 227 177
rect 229 175 234 177
rect 102 163 104 166
rect 75 157 77 162
rect 82 157 84 162
rect 102 161 107 163
rect 105 153 107 161
rect 118 157 120 161
rect 128 153 130 161
rect 176 160 178 164
rect 225 173 234 175
rect 250 175 252 178
rect 232 170 234 173
rect 242 170 244 174
rect 250 173 254 175
rect 252 170 254 173
rect 259 170 261 179
rect 287 173 289 186
rect 297 184 299 195
rect 322 202 328 204
rect 322 200 324 202
rect 326 200 328 202
rect 322 198 331 200
rect 329 195 331 198
rect 307 184 309 188
rect 293 182 299 184
rect 293 180 295 182
rect 297 180 299 182
rect 293 178 299 180
rect 303 182 309 184
rect 303 180 305 182
rect 307 180 309 182
rect 303 178 309 180
rect 294 173 296 178
rect 307 173 309 178
rect 216 163 218 166
rect 138 153 140 158
rect 145 153 147 158
rect 105 151 130 153
rect 189 157 191 162
rect 196 157 198 162
rect 216 161 221 163
rect 219 153 221 161
rect 232 157 234 161
rect 242 153 244 161
rect 329 169 331 187
rect 339 184 341 199
rect 346 194 348 199
rect 345 192 351 194
rect 345 190 347 192
rect 349 190 351 192
rect 345 188 351 190
rect 356 184 358 199
rect 363 189 365 199
rect 443 202 449 204
rect 443 200 445 202
rect 447 200 449 202
rect 335 182 341 184
rect 335 180 337 182
rect 339 180 341 182
rect 335 178 341 180
rect 339 169 341 178
rect 346 182 358 184
rect 362 187 368 189
rect 362 185 364 187
rect 366 185 368 187
rect 362 183 368 185
rect 346 169 348 182
rect 352 176 358 178
rect 352 174 354 176
rect 356 174 358 176
rect 352 172 358 174
rect 356 169 358 172
rect 363 169 365 183
rect 373 179 375 197
rect 396 179 398 197
rect 406 189 408 199
rect 403 187 409 189
rect 403 185 405 187
rect 407 185 409 187
rect 403 183 409 185
rect 413 184 415 199
rect 423 194 425 199
rect 420 192 426 194
rect 420 190 422 192
rect 424 190 426 192
rect 420 188 426 190
rect 430 184 432 199
rect 440 198 449 200
rect 440 195 442 198
rect 542 215 544 219
rect 549 215 551 219
rect 571 215 573 219
rect 529 205 531 210
rect 510 202 516 204
rect 510 200 512 202
rect 514 200 516 202
rect 370 177 376 179
rect 370 175 372 177
rect 374 175 376 177
rect 370 173 376 175
rect 395 177 401 179
rect 395 175 397 177
rect 399 175 401 177
rect 395 173 401 175
rect 373 170 375 173
rect 396 170 398 173
rect 252 153 254 158
rect 259 153 261 158
rect 287 157 289 162
rect 294 157 296 162
rect 219 151 244 153
rect 307 160 309 164
rect 329 153 331 163
rect 406 169 408 183
rect 413 182 425 184
rect 413 176 419 178
rect 413 174 415 176
rect 417 174 419 176
rect 413 172 419 174
rect 413 169 415 172
rect 423 169 425 182
rect 430 182 436 184
rect 430 180 432 182
rect 434 180 436 182
rect 430 178 436 180
rect 430 169 432 178
rect 440 169 442 187
rect 463 179 465 197
rect 473 189 475 199
rect 470 187 476 189
rect 470 185 472 187
rect 474 185 476 187
rect 470 183 476 185
rect 480 184 482 199
rect 490 194 492 199
rect 487 192 493 194
rect 487 190 489 192
rect 491 190 493 192
rect 487 188 493 190
rect 497 184 499 199
rect 507 198 516 200
rect 507 195 509 198
rect 462 177 468 179
rect 462 175 464 177
rect 466 175 468 177
rect 462 173 468 175
rect 463 170 465 173
rect 339 157 341 161
rect 346 153 348 161
rect 356 156 358 161
rect 363 156 365 161
rect 373 156 375 161
rect 396 156 398 161
rect 406 156 408 161
rect 413 156 415 161
rect 329 151 348 153
rect 423 153 425 161
rect 430 157 432 161
rect 440 153 442 163
rect 473 169 475 183
rect 480 182 492 184
rect 480 176 486 178
rect 480 174 482 176
rect 484 174 486 176
rect 480 172 486 174
rect 480 169 482 172
rect 490 169 492 182
rect 497 182 503 184
rect 497 180 499 182
rect 501 180 503 182
rect 497 178 503 180
rect 497 169 499 178
rect 507 169 509 187
rect 529 184 531 187
rect 542 184 544 194
rect 549 191 551 194
rect 549 189 555 191
rect 549 187 551 189
rect 553 187 555 189
rect 607 215 609 219
rect 581 206 583 210
rect 591 206 593 210
rect 618 190 624 192
rect 618 188 620 190
rect 622 188 624 190
rect 549 185 555 187
rect 571 185 573 188
rect 529 182 535 184
rect 529 180 531 182
rect 533 180 535 182
rect 529 178 535 180
rect 539 182 545 184
rect 539 180 541 182
rect 543 180 545 182
rect 539 178 545 180
rect 529 175 531 178
rect 539 175 541 178
rect 549 175 551 185
rect 571 183 577 185
rect 571 181 573 183
rect 575 181 577 183
rect 571 179 577 181
rect 581 184 583 188
rect 591 185 593 188
rect 607 185 609 188
rect 618 186 624 188
rect 618 185 620 186
rect 581 182 587 184
rect 591 183 601 185
rect 607 183 620 185
rect 581 180 583 182
rect 585 180 587 182
rect 572 170 574 179
rect 581 178 587 180
rect 599 179 601 183
rect 581 175 583 178
rect 579 173 583 175
rect 599 177 608 179
rect 599 175 604 177
rect 606 175 608 177
rect 615 175 617 183
rect 579 170 581 173
rect 589 170 591 174
rect 599 173 608 175
rect 599 170 601 173
rect 463 156 465 161
rect 473 156 475 161
rect 480 156 482 161
rect 423 151 442 153
rect 490 153 492 161
rect 497 157 499 161
rect 507 153 509 163
rect 529 161 531 166
rect 539 164 541 169
rect 549 164 551 169
rect 490 151 509 153
rect 615 163 617 166
rect 612 161 617 163
rect 572 153 574 158
rect 579 153 581 158
rect 589 153 591 161
rect 599 157 601 161
rect 612 153 614 161
rect 589 151 614 153
rect 13 132 15 137
rect 23 129 25 134
rect 33 129 35 134
rect 62 134 64 138
rect 75 136 77 141
rect 82 136 84 141
rect 105 145 130 147
rect 105 137 107 145
rect 118 137 120 141
rect 128 137 130 145
rect 138 140 140 145
rect 145 140 147 145
rect 102 135 107 137
rect 102 132 104 135
rect 13 120 15 123
rect 23 120 25 123
rect 13 118 19 120
rect 13 116 15 118
rect 17 116 19 118
rect 13 114 19 116
rect 23 118 29 120
rect 23 116 25 118
rect 27 116 29 118
rect 23 114 29 116
rect 13 111 15 114
rect 26 104 28 114
rect 33 113 35 123
rect 62 120 64 125
rect 75 120 77 125
rect 62 118 68 120
rect 62 116 64 118
rect 66 116 68 118
rect 62 114 68 116
rect 72 118 78 120
rect 72 116 74 118
rect 76 116 78 118
rect 72 114 78 116
rect 33 111 39 113
rect 33 109 35 111
rect 37 109 39 111
rect 62 110 64 114
rect 33 107 39 109
rect 33 104 35 107
rect 13 88 15 93
rect 72 103 74 114
rect 82 112 84 125
rect 176 134 178 138
rect 189 136 191 141
rect 196 136 198 141
rect 219 145 244 147
rect 219 137 221 145
rect 232 137 234 141
rect 242 137 244 145
rect 252 140 254 145
rect 259 140 261 145
rect 118 125 120 128
rect 111 123 120 125
rect 128 124 130 128
rect 138 125 140 128
rect 102 115 104 123
rect 111 121 113 123
rect 115 121 120 123
rect 111 119 120 121
rect 136 123 140 125
rect 136 120 138 123
rect 118 115 120 119
rect 132 118 138 120
rect 145 119 147 128
rect 216 135 221 137
rect 216 132 218 135
rect 176 120 178 125
rect 189 120 191 125
rect 132 116 134 118
rect 136 116 138 118
rect 99 113 112 115
rect 118 113 128 115
rect 132 114 138 116
rect 99 112 101 113
rect 82 110 88 112
rect 82 108 84 110
rect 86 108 88 110
rect 82 106 88 108
rect 95 110 101 112
rect 110 110 112 113
rect 126 110 128 113
rect 136 110 138 114
rect 142 117 148 119
rect 142 115 144 117
rect 146 115 148 117
rect 142 113 148 115
rect 146 110 148 113
rect 176 118 182 120
rect 176 116 178 118
rect 180 116 182 118
rect 176 114 182 116
rect 186 118 192 120
rect 186 116 188 118
rect 190 116 192 118
rect 186 114 192 116
rect 176 110 178 114
rect 95 108 97 110
rect 99 108 101 110
rect 95 106 101 108
rect 82 103 84 106
rect 62 88 64 92
rect 72 85 74 90
rect 82 85 84 90
rect 26 79 28 83
rect 33 79 35 83
rect 126 88 128 92
rect 136 88 138 92
rect 110 79 112 83
rect 186 103 188 114
rect 196 112 198 125
rect 287 136 289 141
rect 294 136 296 141
rect 329 145 348 147
rect 232 125 234 128
rect 225 123 234 125
rect 242 124 244 128
rect 252 125 254 128
rect 216 115 218 123
rect 225 121 227 123
rect 229 121 234 123
rect 225 119 234 121
rect 250 123 254 125
rect 250 120 252 123
rect 232 115 234 119
rect 246 118 252 120
rect 259 119 261 128
rect 307 134 309 138
rect 329 135 331 145
rect 339 137 341 141
rect 346 137 348 145
rect 423 145 442 147
rect 356 137 358 142
rect 363 137 365 142
rect 373 137 375 142
rect 396 137 398 142
rect 406 137 408 142
rect 413 137 415 142
rect 423 137 425 145
rect 430 137 432 141
rect 246 116 248 118
rect 250 116 252 118
rect 213 113 226 115
rect 232 113 242 115
rect 246 114 252 116
rect 213 112 215 113
rect 196 110 202 112
rect 196 108 198 110
rect 200 108 202 110
rect 196 106 202 108
rect 209 110 215 112
rect 224 110 226 113
rect 240 110 242 113
rect 250 110 252 114
rect 256 117 262 119
rect 256 115 258 117
rect 260 115 262 117
rect 256 113 262 115
rect 260 110 262 113
rect 287 112 289 125
rect 294 120 296 125
rect 307 120 309 125
rect 293 118 299 120
rect 293 116 295 118
rect 297 116 299 118
rect 293 114 299 116
rect 303 118 309 120
rect 303 116 305 118
rect 307 116 309 118
rect 303 114 309 116
rect 283 110 289 112
rect 209 108 211 110
rect 213 108 215 110
rect 209 106 215 108
rect 196 103 198 106
rect 176 88 178 92
rect 186 85 188 90
rect 196 85 198 90
rect 146 79 148 83
rect 240 88 242 92
rect 250 88 252 92
rect 224 79 226 83
rect 283 108 285 110
rect 287 108 289 110
rect 283 106 289 108
rect 287 103 289 106
rect 297 103 299 114
rect 307 110 309 114
rect 329 111 331 129
rect 339 120 341 129
rect 335 118 341 120
rect 335 116 337 118
rect 339 116 341 118
rect 335 114 341 116
rect 346 116 348 129
rect 356 126 358 129
rect 352 124 358 126
rect 352 122 354 124
rect 356 122 358 124
rect 352 120 358 122
rect 346 114 358 116
rect 363 115 365 129
rect 440 135 442 145
rect 490 145 509 147
rect 463 137 465 142
rect 473 137 475 142
rect 480 137 482 142
rect 490 137 492 145
rect 497 137 499 141
rect 373 125 375 128
rect 396 125 398 128
rect 370 123 376 125
rect 370 121 372 123
rect 374 121 376 123
rect 370 119 376 121
rect 395 123 401 125
rect 395 121 397 123
rect 399 121 401 123
rect 395 119 401 121
rect 329 100 331 103
rect 322 98 331 100
rect 339 99 341 114
rect 345 108 351 110
rect 345 106 347 108
rect 349 106 351 108
rect 345 104 351 106
rect 346 99 348 104
rect 356 99 358 114
rect 362 113 368 115
rect 362 111 364 113
rect 366 111 368 113
rect 362 109 368 111
rect 363 99 365 109
rect 373 101 375 119
rect 396 101 398 119
rect 406 115 408 129
rect 413 126 415 129
rect 413 124 419 126
rect 413 122 415 124
rect 417 122 419 124
rect 413 120 419 122
rect 423 116 425 129
rect 403 113 409 115
rect 403 111 405 113
rect 407 111 409 113
rect 403 109 409 111
rect 413 114 425 116
rect 430 120 432 129
rect 430 118 436 120
rect 430 116 432 118
rect 434 116 436 118
rect 430 114 436 116
rect 322 96 324 98
rect 326 96 328 98
rect 322 94 328 96
rect 287 85 289 90
rect 297 85 299 90
rect 307 88 309 92
rect 260 79 262 83
rect 406 99 408 109
rect 413 99 415 114
rect 420 108 426 110
rect 420 106 422 108
rect 424 106 426 108
rect 420 104 426 106
rect 423 99 425 104
rect 430 99 432 114
rect 440 111 442 129
rect 507 135 509 145
rect 589 145 614 147
rect 529 132 531 137
rect 463 125 465 128
rect 462 123 468 125
rect 462 121 464 123
rect 466 121 468 123
rect 462 119 468 121
rect 440 100 442 103
rect 463 101 465 119
rect 473 115 475 129
rect 480 126 482 129
rect 480 124 486 126
rect 480 122 482 124
rect 484 122 486 124
rect 480 120 486 122
rect 490 116 492 129
rect 470 113 476 115
rect 470 111 472 113
rect 474 111 476 113
rect 470 109 476 111
rect 480 114 492 116
rect 497 120 499 129
rect 497 118 503 120
rect 497 116 499 118
rect 501 116 503 118
rect 497 114 503 116
rect 440 98 449 100
rect 443 96 445 98
rect 447 96 449 98
rect 443 94 449 96
rect 473 99 475 109
rect 480 99 482 114
rect 487 108 493 110
rect 487 106 489 108
rect 491 106 493 108
rect 487 104 493 106
rect 490 99 492 104
rect 497 99 499 114
rect 507 111 509 129
rect 539 129 541 134
rect 549 129 551 134
rect 572 140 574 145
rect 579 140 581 145
rect 589 137 591 145
rect 599 137 601 141
rect 612 137 614 145
rect 612 135 617 137
rect 615 132 617 135
rect 529 120 531 123
rect 539 120 541 123
rect 529 118 535 120
rect 529 116 531 118
rect 533 116 535 118
rect 529 114 535 116
rect 539 118 545 120
rect 539 116 541 118
rect 543 116 545 118
rect 539 114 545 116
rect 529 111 531 114
rect 507 100 509 103
rect 507 98 516 100
rect 510 96 512 98
rect 514 96 516 98
rect 510 94 516 96
rect 542 104 544 114
rect 549 113 551 123
rect 572 119 574 128
rect 579 125 581 128
rect 579 123 583 125
rect 589 124 591 128
rect 599 125 601 128
rect 581 120 583 123
rect 599 123 608 125
rect 599 121 604 123
rect 606 121 608 123
rect 571 117 577 119
rect 571 115 573 117
rect 575 115 577 117
rect 571 113 577 115
rect 581 118 587 120
rect 581 116 583 118
rect 585 116 587 118
rect 581 114 587 116
rect 599 119 608 121
rect 599 115 601 119
rect 615 115 617 123
rect 549 111 555 113
rect 549 109 551 111
rect 553 109 555 111
rect 571 110 573 113
rect 581 110 583 114
rect 591 113 601 115
rect 607 113 620 115
rect 591 110 593 113
rect 607 110 609 113
rect 618 112 620 113
rect 618 110 624 112
rect 549 107 555 109
rect 549 104 551 107
rect 529 88 531 93
rect 339 79 341 83
rect 346 79 348 83
rect 356 79 358 83
rect 363 79 365 83
rect 373 79 375 83
rect 396 79 398 83
rect 406 79 408 83
rect 413 79 415 83
rect 423 79 425 83
rect 430 79 432 83
rect 463 79 465 83
rect 473 79 475 83
rect 480 79 482 83
rect 490 79 492 83
rect 497 79 499 83
rect 581 88 583 92
rect 591 88 593 92
rect 542 79 544 83
rect 549 79 551 83
rect 571 79 573 83
rect 618 108 620 110
rect 622 108 624 110
rect 618 106 624 108
rect 607 79 609 83
rect 26 71 28 75
rect 33 71 35 75
rect 13 61 15 66
rect 110 71 112 75
rect 62 62 64 66
rect 72 64 74 69
rect 82 64 84 69
rect 13 40 15 43
rect 26 40 28 50
rect 33 47 35 50
rect 33 45 39 47
rect 33 43 35 45
rect 37 43 39 45
rect 33 41 39 43
rect 13 38 19 40
rect 13 36 15 38
rect 17 36 19 38
rect 13 34 19 36
rect 23 38 29 40
rect 23 36 25 38
rect 27 36 29 38
rect 23 34 29 36
rect 13 31 15 34
rect 23 31 25 34
rect 33 31 35 41
rect 62 40 64 44
rect 72 40 74 51
rect 82 48 84 51
rect 82 46 88 48
rect 82 44 84 46
rect 86 44 88 46
rect 82 42 88 44
rect 95 46 101 48
rect 95 44 97 46
rect 99 44 101 46
rect 146 71 148 75
rect 126 62 128 66
rect 136 62 138 66
rect 224 71 226 75
rect 176 62 178 66
rect 186 64 188 69
rect 196 64 198 69
rect 95 42 101 44
rect 62 38 68 40
rect 62 36 64 38
rect 66 36 68 38
rect 62 34 68 36
rect 72 38 78 40
rect 72 36 74 38
rect 76 36 78 38
rect 72 34 78 36
rect 62 29 64 34
rect 75 29 77 34
rect 82 29 84 42
rect 99 41 101 42
rect 110 41 112 44
rect 126 41 128 44
rect 99 39 112 41
rect 118 39 128 41
rect 136 40 138 44
rect 146 41 148 44
rect 102 31 104 39
rect 118 35 120 39
rect 111 33 120 35
rect 132 38 138 40
rect 132 36 134 38
rect 136 36 138 38
rect 132 34 138 36
rect 142 39 148 41
rect 142 37 144 39
rect 146 37 148 39
rect 142 35 148 37
rect 176 40 178 44
rect 186 40 188 51
rect 196 48 198 51
rect 196 46 202 48
rect 196 44 198 46
rect 200 44 202 46
rect 196 42 202 44
rect 209 46 215 48
rect 209 44 211 46
rect 213 44 215 46
rect 260 71 262 75
rect 240 62 242 66
rect 250 62 252 66
rect 339 71 341 75
rect 346 71 348 75
rect 356 71 358 75
rect 363 71 365 75
rect 373 71 375 75
rect 396 71 398 75
rect 406 71 408 75
rect 413 71 415 75
rect 423 71 425 75
rect 430 71 432 75
rect 463 71 465 75
rect 473 71 475 75
rect 480 71 482 75
rect 490 71 492 75
rect 497 71 499 75
rect 287 64 289 69
rect 297 64 299 69
rect 307 62 309 66
rect 287 48 289 51
rect 283 46 289 48
rect 283 44 285 46
rect 287 44 289 46
rect 209 42 215 44
rect 176 38 182 40
rect 176 36 178 38
rect 180 36 182 38
rect 111 31 113 33
rect 115 31 120 33
rect 13 17 15 22
rect 23 20 25 25
rect 33 20 35 25
rect 62 16 64 20
rect 111 29 120 31
rect 136 31 138 34
rect 118 26 120 29
rect 128 26 130 30
rect 136 29 140 31
rect 138 26 140 29
rect 145 26 147 35
rect 176 34 182 36
rect 186 38 192 40
rect 186 36 188 38
rect 190 36 192 38
rect 186 34 192 36
rect 176 29 178 34
rect 189 29 191 34
rect 196 29 198 42
rect 213 41 215 42
rect 224 41 226 44
rect 240 41 242 44
rect 213 39 226 41
rect 232 39 242 41
rect 250 40 252 44
rect 260 41 262 44
rect 283 42 289 44
rect 216 31 218 39
rect 232 35 234 39
rect 225 33 234 35
rect 246 38 252 40
rect 246 36 248 38
rect 250 36 252 38
rect 246 34 252 36
rect 256 39 262 41
rect 256 37 258 39
rect 260 37 262 39
rect 256 35 262 37
rect 225 31 227 33
rect 229 31 234 33
rect 102 19 104 22
rect 75 13 77 18
rect 82 13 84 18
rect 102 17 107 19
rect 105 9 107 17
rect 118 13 120 17
rect 128 9 130 17
rect 176 16 178 20
rect 225 29 234 31
rect 250 31 252 34
rect 232 26 234 29
rect 242 26 244 30
rect 250 29 254 31
rect 252 26 254 29
rect 259 26 261 35
rect 287 29 289 42
rect 297 40 299 51
rect 322 58 328 60
rect 322 56 324 58
rect 326 56 328 58
rect 322 54 331 56
rect 329 51 331 54
rect 307 40 309 44
rect 293 38 299 40
rect 293 36 295 38
rect 297 36 299 38
rect 293 34 299 36
rect 303 38 309 40
rect 303 36 305 38
rect 307 36 309 38
rect 303 34 309 36
rect 294 29 296 34
rect 307 29 309 34
rect 216 19 218 22
rect 138 9 140 14
rect 145 9 147 14
rect 105 7 130 9
rect 189 13 191 18
rect 196 13 198 18
rect 216 17 221 19
rect 219 9 221 17
rect 232 13 234 17
rect 242 9 244 17
rect 329 25 331 43
rect 339 40 341 55
rect 346 50 348 55
rect 345 48 351 50
rect 345 46 347 48
rect 349 46 351 48
rect 345 44 351 46
rect 356 40 358 55
rect 363 45 365 55
rect 443 58 449 60
rect 443 56 445 58
rect 447 56 449 58
rect 335 38 341 40
rect 335 36 337 38
rect 339 36 341 38
rect 335 34 341 36
rect 339 25 341 34
rect 346 38 358 40
rect 362 43 368 45
rect 362 41 364 43
rect 366 41 368 43
rect 362 39 368 41
rect 346 25 348 38
rect 352 32 358 34
rect 352 30 354 32
rect 356 30 358 32
rect 352 28 358 30
rect 356 25 358 28
rect 363 25 365 39
rect 373 35 375 53
rect 396 35 398 53
rect 406 45 408 55
rect 403 43 409 45
rect 403 41 405 43
rect 407 41 409 43
rect 403 39 409 41
rect 413 40 415 55
rect 423 50 425 55
rect 420 48 426 50
rect 420 46 422 48
rect 424 46 426 48
rect 420 44 426 46
rect 430 40 432 55
rect 440 54 449 56
rect 440 51 442 54
rect 542 71 544 75
rect 549 71 551 75
rect 571 71 573 75
rect 529 61 531 66
rect 510 58 516 60
rect 510 56 512 58
rect 514 56 516 58
rect 370 33 376 35
rect 370 31 372 33
rect 374 31 376 33
rect 370 29 376 31
rect 395 33 401 35
rect 395 31 397 33
rect 399 31 401 33
rect 395 29 401 31
rect 373 26 375 29
rect 396 26 398 29
rect 252 9 254 14
rect 259 9 261 14
rect 287 13 289 18
rect 294 13 296 18
rect 219 7 244 9
rect 307 16 309 20
rect 329 9 331 19
rect 406 25 408 39
rect 413 38 425 40
rect 413 32 419 34
rect 413 30 415 32
rect 417 30 419 32
rect 413 28 419 30
rect 413 25 415 28
rect 423 25 425 38
rect 430 38 436 40
rect 430 36 432 38
rect 434 36 436 38
rect 430 34 436 36
rect 430 25 432 34
rect 440 25 442 43
rect 463 35 465 53
rect 473 45 475 55
rect 470 43 476 45
rect 470 41 472 43
rect 474 41 476 43
rect 470 39 476 41
rect 480 40 482 55
rect 490 50 492 55
rect 487 48 493 50
rect 487 46 489 48
rect 491 46 493 48
rect 487 44 493 46
rect 497 40 499 55
rect 507 54 516 56
rect 507 51 509 54
rect 462 33 468 35
rect 462 31 464 33
rect 466 31 468 33
rect 462 29 468 31
rect 463 26 465 29
rect 339 13 341 17
rect 346 9 348 17
rect 356 12 358 17
rect 363 12 365 17
rect 373 12 375 17
rect 396 12 398 17
rect 406 12 408 17
rect 413 12 415 17
rect 329 7 348 9
rect 423 9 425 17
rect 430 13 432 17
rect 440 9 442 19
rect 473 25 475 39
rect 480 38 492 40
rect 480 32 486 34
rect 480 30 482 32
rect 484 30 486 32
rect 480 28 486 30
rect 480 25 482 28
rect 490 25 492 38
rect 497 38 503 40
rect 497 36 499 38
rect 501 36 503 38
rect 497 34 503 36
rect 497 25 499 34
rect 507 25 509 43
rect 529 40 531 43
rect 542 40 544 50
rect 549 47 551 50
rect 549 45 555 47
rect 549 43 551 45
rect 553 43 555 45
rect 607 71 609 75
rect 581 62 583 66
rect 591 62 593 66
rect 618 46 624 48
rect 618 44 620 46
rect 622 44 624 46
rect 549 41 555 43
rect 571 41 573 44
rect 529 38 535 40
rect 529 36 531 38
rect 533 36 535 38
rect 529 34 535 36
rect 539 38 545 40
rect 539 36 541 38
rect 543 36 545 38
rect 539 34 545 36
rect 529 31 531 34
rect 539 31 541 34
rect 549 31 551 41
rect 571 39 577 41
rect 571 37 573 39
rect 575 37 577 39
rect 571 35 577 37
rect 581 40 583 44
rect 591 41 593 44
rect 607 41 609 44
rect 618 42 624 44
rect 618 41 620 42
rect 581 38 587 40
rect 591 39 601 41
rect 607 39 620 41
rect 581 36 583 38
rect 585 36 587 38
rect 572 26 574 35
rect 581 34 587 36
rect 599 35 601 39
rect 581 31 583 34
rect 579 29 583 31
rect 599 33 608 35
rect 599 31 604 33
rect 606 31 608 33
rect 615 31 617 39
rect 579 26 581 29
rect 589 26 591 30
rect 599 29 608 31
rect 599 26 601 29
rect 463 12 465 17
rect 473 12 475 17
rect 480 12 482 17
rect 423 7 442 9
rect 490 9 492 17
rect 497 13 499 17
rect 507 9 509 19
rect 529 17 531 22
rect 539 20 541 25
rect 549 20 551 25
rect 490 7 509 9
rect 615 19 617 22
rect 612 17 617 19
rect 572 9 574 14
rect 579 9 581 14
rect 589 9 591 17
rect 599 13 601 17
rect 612 9 614 17
rect 589 7 614 9
<< ndif >>
rect 17 572 23 574
rect 17 570 19 572
rect 21 570 23 572
rect 17 568 23 570
rect 36 572 42 574
rect 66 576 73 578
rect 66 574 68 576
rect 70 574 73 576
rect 36 570 38 572
rect 40 570 42 572
rect 36 568 42 570
rect 17 564 21 568
rect 8 561 13 564
rect 6 559 13 561
rect 6 557 8 559
rect 10 557 13 559
rect 6 555 13 557
rect 15 561 21 564
rect 37 561 42 568
rect 66 568 73 574
rect 149 576 155 578
rect 149 574 151 576
rect 153 574 155 576
rect 149 572 155 574
rect 180 576 187 578
rect 180 574 182 576
rect 184 574 187 576
rect 133 569 138 572
rect 66 566 75 568
rect 15 555 23 561
rect 25 559 33 561
rect 25 557 28 559
rect 30 557 33 559
rect 25 555 33 557
rect 35 555 42 561
rect 55 564 62 566
rect 55 562 57 564
rect 59 562 62 564
rect 55 560 62 562
rect 57 557 62 560
rect 64 557 75 566
rect 77 557 82 568
rect 84 566 91 568
rect 84 564 87 566
rect 89 564 91 566
rect 109 567 118 569
rect 109 565 111 567
rect 113 565 118 567
rect 109 564 118 565
rect 84 562 91 564
rect 84 557 89 562
rect 97 561 102 564
rect 95 559 102 561
rect 95 557 97 559
rect 99 557 102 559
rect 95 555 102 557
rect 104 560 118 564
rect 120 564 128 569
rect 120 562 123 564
rect 125 562 128 564
rect 120 560 128 562
rect 130 566 138 569
rect 130 564 133 566
rect 135 564 138 566
rect 130 560 138 564
rect 140 560 145 572
rect 147 560 155 572
rect 180 568 187 574
rect 263 576 269 578
rect 263 574 265 576
rect 267 574 269 576
rect 263 572 269 574
rect 298 576 305 578
rect 298 574 301 576
rect 303 574 305 576
rect 247 569 252 572
rect 180 566 189 568
rect 169 564 176 566
rect 169 562 171 564
rect 173 562 176 564
rect 169 560 176 562
rect 104 555 109 560
rect 171 557 176 560
rect 178 557 189 566
rect 191 557 196 568
rect 198 566 205 568
rect 198 564 201 566
rect 203 564 205 566
rect 223 567 232 569
rect 223 565 225 567
rect 227 565 232 567
rect 223 564 232 565
rect 198 562 205 564
rect 198 557 203 562
rect 211 561 216 564
rect 209 559 216 561
rect 209 557 211 559
rect 213 557 216 559
rect 209 555 216 557
rect 218 560 232 564
rect 234 564 242 569
rect 234 562 237 564
rect 239 562 242 564
rect 234 560 242 562
rect 244 566 252 569
rect 244 564 247 566
rect 249 564 252 566
rect 244 560 252 564
rect 254 560 259 572
rect 261 560 269 572
rect 298 568 305 574
rect 280 566 287 568
rect 280 564 282 566
rect 284 564 287 566
rect 280 562 287 564
rect 218 555 223 560
rect 282 557 287 562
rect 289 557 294 568
rect 296 566 305 568
rect 333 567 339 569
rect 296 557 307 566
rect 309 564 316 566
rect 309 562 312 564
rect 314 562 316 564
rect 309 560 316 562
rect 322 565 329 567
rect 322 563 324 565
rect 326 563 329 565
rect 322 561 329 563
rect 331 565 339 567
rect 331 563 334 565
rect 336 563 339 565
rect 331 561 339 563
rect 341 561 346 569
rect 348 567 356 569
rect 348 565 351 567
rect 353 565 356 567
rect 348 561 356 565
rect 358 561 363 569
rect 365 567 373 569
rect 365 565 368 567
rect 370 565 373 567
rect 365 561 373 565
rect 309 557 314 560
rect 368 560 373 561
rect 375 566 380 569
rect 391 566 396 569
rect 375 564 382 566
rect 375 562 378 564
rect 380 562 382 564
rect 375 560 382 562
rect 389 564 396 566
rect 389 562 391 564
rect 393 562 396 564
rect 389 560 396 562
rect 398 567 406 569
rect 398 565 401 567
rect 403 565 406 567
rect 398 561 406 565
rect 408 561 413 569
rect 415 567 423 569
rect 415 565 418 567
rect 420 565 423 567
rect 415 561 423 565
rect 425 561 430 569
rect 432 567 438 569
rect 432 565 440 567
rect 432 563 435 565
rect 437 563 440 565
rect 432 561 440 563
rect 442 565 449 567
rect 458 566 463 569
rect 442 563 445 565
rect 447 563 449 565
rect 442 561 449 563
rect 456 564 463 566
rect 456 562 458 564
rect 460 562 463 564
rect 398 560 403 561
rect 456 560 463 562
rect 465 567 473 569
rect 465 565 468 567
rect 470 565 473 567
rect 465 561 473 565
rect 475 561 480 569
rect 482 567 490 569
rect 482 565 485 567
rect 487 565 490 567
rect 482 561 490 565
rect 492 561 497 569
rect 499 567 505 569
rect 564 576 570 578
rect 564 574 566 576
rect 568 574 570 576
rect 533 572 539 574
rect 533 570 535 572
rect 537 570 539 572
rect 499 565 507 567
rect 499 563 502 565
rect 504 563 507 565
rect 499 561 507 563
rect 509 565 516 567
rect 509 563 512 565
rect 514 563 516 565
rect 533 568 539 570
rect 552 572 558 574
rect 552 570 554 572
rect 556 570 558 572
rect 552 568 558 570
rect 533 564 537 568
rect 509 561 516 563
rect 524 561 529 564
rect 465 560 470 561
rect 522 559 529 561
rect 522 557 524 559
rect 526 557 529 559
rect 522 555 529 557
rect 531 561 537 564
rect 553 561 558 568
rect 531 555 539 561
rect 541 559 549 561
rect 541 557 544 559
rect 546 557 549 559
rect 541 555 549 557
rect 551 555 558 561
rect 564 572 570 574
rect 564 560 572 572
rect 574 560 579 572
rect 581 569 586 572
rect 581 566 589 569
rect 581 564 584 566
rect 586 564 589 566
rect 581 560 589 564
rect 591 564 599 569
rect 591 562 594 564
rect 596 562 599 564
rect 591 560 599 562
rect 601 567 610 569
rect 601 565 606 567
rect 608 565 610 567
rect 601 564 610 565
rect 601 560 615 564
rect 610 555 615 560
rect 617 561 622 564
rect 617 559 624 561
rect 617 557 620 559
rect 622 557 624 559
rect 617 555 624 557
rect 6 461 13 463
rect 6 459 8 461
rect 10 459 13 461
rect 6 457 13 459
rect 8 454 13 457
rect 15 457 23 463
rect 25 461 33 463
rect 25 459 28 461
rect 30 459 33 461
rect 25 457 33 459
rect 35 457 42 463
rect 95 461 102 463
rect 57 458 62 461
rect 15 454 21 457
rect 17 450 21 454
rect 37 450 42 457
rect 55 456 62 458
rect 55 454 57 456
rect 59 454 62 456
rect 55 452 62 454
rect 64 452 75 461
rect 17 448 23 450
rect 17 446 19 448
rect 21 446 23 448
rect 17 444 23 446
rect 36 448 42 450
rect 66 450 75 452
rect 77 450 82 461
rect 84 456 89 461
rect 95 459 97 461
rect 99 459 102 461
rect 95 457 102 459
rect 84 454 91 456
rect 97 454 102 457
rect 104 458 109 463
rect 209 461 216 463
rect 171 458 176 461
rect 104 454 118 458
rect 84 452 87 454
rect 89 452 91 454
rect 84 450 91 452
rect 109 453 118 454
rect 109 451 111 453
rect 113 451 118 453
rect 36 446 38 448
rect 40 446 42 448
rect 36 444 42 446
rect 66 444 73 450
rect 109 449 118 451
rect 120 456 128 458
rect 120 454 123 456
rect 125 454 128 456
rect 120 449 128 454
rect 130 454 138 458
rect 130 452 133 454
rect 135 452 138 454
rect 130 449 138 452
rect 66 442 68 444
rect 70 442 73 444
rect 66 440 73 442
rect 133 446 138 449
rect 140 446 145 458
rect 147 446 155 458
rect 169 456 176 458
rect 169 454 171 456
rect 173 454 176 456
rect 169 452 176 454
rect 178 452 189 461
rect 180 450 189 452
rect 191 450 196 461
rect 198 456 203 461
rect 209 459 211 461
rect 213 459 216 461
rect 209 457 216 459
rect 198 454 205 456
rect 211 454 216 457
rect 218 458 223 463
rect 218 454 232 458
rect 198 452 201 454
rect 203 452 205 454
rect 198 450 205 452
rect 223 453 232 454
rect 223 451 225 453
rect 227 451 232 453
rect 149 444 155 446
rect 149 442 151 444
rect 153 442 155 444
rect 149 440 155 442
rect 180 444 187 450
rect 223 449 232 451
rect 234 456 242 458
rect 234 454 237 456
rect 239 454 242 456
rect 234 449 242 454
rect 244 454 252 458
rect 244 452 247 454
rect 249 452 252 454
rect 244 449 252 452
rect 180 442 182 444
rect 184 442 187 444
rect 180 440 187 442
rect 247 446 252 449
rect 254 446 259 458
rect 261 446 269 458
rect 282 456 287 461
rect 280 454 287 456
rect 280 452 282 454
rect 284 452 287 454
rect 280 450 287 452
rect 289 450 294 461
rect 296 452 307 461
rect 309 458 314 461
rect 309 456 316 458
rect 368 457 373 458
rect 309 454 312 456
rect 314 454 316 456
rect 309 452 316 454
rect 322 455 329 457
rect 322 453 324 455
rect 326 453 329 455
rect 296 450 305 452
rect 263 444 269 446
rect 263 442 265 444
rect 267 442 269 444
rect 263 440 269 442
rect 298 444 305 450
rect 322 451 329 453
rect 331 455 339 457
rect 331 453 334 455
rect 336 453 339 455
rect 331 451 339 453
rect 298 442 301 444
rect 303 442 305 444
rect 298 440 305 442
rect 333 449 339 451
rect 341 449 346 457
rect 348 453 356 457
rect 348 451 351 453
rect 353 451 356 453
rect 348 449 356 451
rect 358 449 363 457
rect 365 453 373 457
rect 365 451 368 453
rect 370 451 373 453
rect 365 449 373 451
rect 375 456 382 458
rect 375 454 378 456
rect 380 454 382 456
rect 375 452 382 454
rect 389 456 396 458
rect 389 454 391 456
rect 393 454 396 456
rect 389 452 396 454
rect 375 449 380 452
rect 391 449 396 452
rect 398 457 403 458
rect 398 453 406 457
rect 398 451 401 453
rect 403 451 406 453
rect 398 449 406 451
rect 408 449 413 457
rect 415 453 423 457
rect 415 451 418 453
rect 420 451 423 453
rect 415 449 423 451
rect 425 449 430 457
rect 432 455 440 457
rect 432 453 435 455
rect 437 453 440 455
rect 432 451 440 453
rect 442 455 449 457
rect 442 453 445 455
rect 447 453 449 455
rect 442 451 449 453
rect 456 456 463 458
rect 456 454 458 456
rect 460 454 463 456
rect 456 452 463 454
rect 432 449 438 451
rect 458 449 463 452
rect 465 457 470 458
rect 522 461 529 463
rect 522 459 524 461
rect 526 459 529 461
rect 522 457 529 459
rect 465 453 473 457
rect 465 451 468 453
rect 470 451 473 453
rect 465 449 473 451
rect 475 449 480 457
rect 482 453 490 457
rect 482 451 485 453
rect 487 451 490 453
rect 482 449 490 451
rect 492 449 497 457
rect 499 455 507 457
rect 499 453 502 455
rect 504 453 507 455
rect 499 451 507 453
rect 509 455 516 457
rect 509 453 512 455
rect 514 453 516 455
rect 524 454 529 457
rect 531 457 539 463
rect 541 461 549 463
rect 541 459 544 461
rect 546 459 549 461
rect 541 457 549 459
rect 551 457 558 463
rect 610 458 615 463
rect 531 454 537 457
rect 509 451 516 453
rect 499 449 505 451
rect 533 450 537 454
rect 553 450 558 457
rect 533 448 539 450
rect 533 446 535 448
rect 537 446 539 448
rect 533 444 539 446
rect 552 448 558 450
rect 552 446 554 448
rect 556 446 558 448
rect 552 444 558 446
rect 564 446 572 458
rect 574 446 579 458
rect 581 454 589 458
rect 581 452 584 454
rect 586 452 589 454
rect 581 449 589 452
rect 591 456 599 458
rect 591 454 594 456
rect 596 454 599 456
rect 591 449 599 454
rect 601 454 615 458
rect 617 461 624 463
rect 617 459 620 461
rect 622 459 624 461
rect 617 457 624 459
rect 617 454 622 457
rect 601 453 610 454
rect 601 451 606 453
rect 608 451 610 453
rect 601 449 610 451
rect 581 446 586 449
rect 564 444 570 446
rect 564 442 566 444
rect 568 442 570 444
rect 564 440 570 442
rect 17 428 23 430
rect 17 426 19 428
rect 21 426 23 428
rect 17 424 23 426
rect 36 428 42 430
rect 66 432 73 434
rect 66 430 68 432
rect 70 430 73 432
rect 36 426 38 428
rect 40 426 42 428
rect 36 424 42 426
rect 17 420 21 424
rect 8 417 13 420
rect 6 415 13 417
rect 6 413 8 415
rect 10 413 13 415
rect 6 411 13 413
rect 15 417 21 420
rect 37 417 42 424
rect 66 424 73 430
rect 149 432 155 434
rect 149 430 151 432
rect 153 430 155 432
rect 149 428 155 430
rect 180 432 187 434
rect 180 430 182 432
rect 184 430 187 432
rect 133 425 138 428
rect 66 422 75 424
rect 15 411 23 417
rect 25 415 33 417
rect 25 413 28 415
rect 30 413 33 415
rect 25 411 33 413
rect 35 411 42 417
rect 55 420 62 422
rect 55 418 57 420
rect 59 418 62 420
rect 55 416 62 418
rect 57 413 62 416
rect 64 413 75 422
rect 77 413 82 424
rect 84 422 91 424
rect 84 420 87 422
rect 89 420 91 422
rect 109 423 118 425
rect 109 421 111 423
rect 113 421 118 423
rect 109 420 118 421
rect 84 418 91 420
rect 84 413 89 418
rect 97 417 102 420
rect 95 415 102 417
rect 95 413 97 415
rect 99 413 102 415
rect 95 411 102 413
rect 104 416 118 420
rect 120 420 128 425
rect 120 418 123 420
rect 125 418 128 420
rect 120 416 128 418
rect 130 422 138 425
rect 130 420 133 422
rect 135 420 138 422
rect 130 416 138 420
rect 140 416 145 428
rect 147 416 155 428
rect 180 424 187 430
rect 263 432 269 434
rect 263 430 265 432
rect 267 430 269 432
rect 263 428 269 430
rect 298 432 305 434
rect 298 430 301 432
rect 303 430 305 432
rect 247 425 252 428
rect 180 422 189 424
rect 169 420 176 422
rect 169 418 171 420
rect 173 418 176 420
rect 169 416 176 418
rect 104 411 109 416
rect 171 413 176 416
rect 178 413 189 422
rect 191 413 196 424
rect 198 422 205 424
rect 198 420 201 422
rect 203 420 205 422
rect 223 423 232 425
rect 223 421 225 423
rect 227 421 232 423
rect 223 420 232 421
rect 198 418 205 420
rect 198 413 203 418
rect 211 417 216 420
rect 209 415 216 417
rect 209 413 211 415
rect 213 413 216 415
rect 209 411 216 413
rect 218 416 232 420
rect 234 420 242 425
rect 234 418 237 420
rect 239 418 242 420
rect 234 416 242 418
rect 244 422 252 425
rect 244 420 247 422
rect 249 420 252 422
rect 244 416 252 420
rect 254 416 259 428
rect 261 416 269 428
rect 298 424 305 430
rect 280 422 287 424
rect 280 420 282 422
rect 284 420 287 422
rect 280 418 287 420
rect 218 411 223 416
rect 282 413 287 418
rect 289 413 294 424
rect 296 422 305 424
rect 333 423 339 425
rect 296 413 307 422
rect 309 420 316 422
rect 309 418 312 420
rect 314 418 316 420
rect 309 416 316 418
rect 322 421 329 423
rect 322 419 324 421
rect 326 419 329 421
rect 322 417 329 419
rect 331 421 339 423
rect 331 419 334 421
rect 336 419 339 421
rect 331 417 339 419
rect 341 417 346 425
rect 348 423 356 425
rect 348 421 351 423
rect 353 421 356 423
rect 348 417 356 421
rect 358 417 363 425
rect 365 423 373 425
rect 365 421 368 423
rect 370 421 373 423
rect 365 417 373 421
rect 309 413 314 416
rect 368 416 373 417
rect 375 422 380 425
rect 391 422 396 425
rect 375 420 382 422
rect 375 418 378 420
rect 380 418 382 420
rect 375 416 382 418
rect 389 420 396 422
rect 389 418 391 420
rect 393 418 396 420
rect 389 416 396 418
rect 398 423 406 425
rect 398 421 401 423
rect 403 421 406 423
rect 398 417 406 421
rect 408 417 413 425
rect 415 423 423 425
rect 415 421 418 423
rect 420 421 423 423
rect 415 417 423 421
rect 425 417 430 425
rect 432 423 438 425
rect 432 421 440 423
rect 432 419 435 421
rect 437 419 440 421
rect 432 417 440 419
rect 442 421 449 423
rect 458 422 463 425
rect 442 419 445 421
rect 447 419 449 421
rect 442 417 449 419
rect 456 420 463 422
rect 456 418 458 420
rect 460 418 463 420
rect 398 416 403 417
rect 456 416 463 418
rect 465 423 473 425
rect 465 421 468 423
rect 470 421 473 423
rect 465 417 473 421
rect 475 417 480 425
rect 482 423 490 425
rect 482 421 485 423
rect 487 421 490 423
rect 482 417 490 421
rect 492 417 497 425
rect 499 423 505 425
rect 564 432 570 434
rect 564 430 566 432
rect 568 430 570 432
rect 533 428 539 430
rect 533 426 535 428
rect 537 426 539 428
rect 499 421 507 423
rect 499 419 502 421
rect 504 419 507 421
rect 499 417 507 419
rect 509 421 516 423
rect 509 419 512 421
rect 514 419 516 421
rect 533 424 539 426
rect 552 428 558 430
rect 552 426 554 428
rect 556 426 558 428
rect 552 424 558 426
rect 533 420 537 424
rect 509 417 516 419
rect 524 417 529 420
rect 465 416 470 417
rect 522 415 529 417
rect 522 413 524 415
rect 526 413 529 415
rect 522 411 529 413
rect 531 417 537 420
rect 553 417 558 424
rect 531 411 539 417
rect 541 415 549 417
rect 541 413 544 415
rect 546 413 549 415
rect 541 411 549 413
rect 551 411 558 417
rect 564 428 570 430
rect 564 416 572 428
rect 574 416 579 428
rect 581 425 586 428
rect 581 422 589 425
rect 581 420 584 422
rect 586 420 589 422
rect 581 416 589 420
rect 591 420 599 425
rect 591 418 594 420
rect 596 418 599 420
rect 591 416 599 418
rect 601 423 610 425
rect 601 421 606 423
rect 608 421 610 423
rect 601 420 610 421
rect 601 416 615 420
rect 610 411 615 416
rect 617 417 622 420
rect 617 415 624 417
rect 617 413 620 415
rect 622 413 624 415
rect 617 411 624 413
rect 6 317 13 319
rect 6 315 8 317
rect 10 315 13 317
rect 6 313 13 315
rect 8 310 13 313
rect 15 313 23 319
rect 25 317 33 319
rect 25 315 28 317
rect 30 315 33 317
rect 25 313 33 315
rect 35 313 42 319
rect 95 317 102 319
rect 57 314 62 317
rect 15 310 21 313
rect 17 306 21 310
rect 37 306 42 313
rect 55 312 62 314
rect 55 310 57 312
rect 59 310 62 312
rect 55 308 62 310
rect 64 308 75 317
rect 17 304 23 306
rect 17 302 19 304
rect 21 302 23 304
rect 17 300 23 302
rect 36 304 42 306
rect 66 306 75 308
rect 77 306 82 317
rect 84 312 89 317
rect 95 315 97 317
rect 99 315 102 317
rect 95 313 102 315
rect 84 310 91 312
rect 97 310 102 313
rect 104 314 109 319
rect 209 317 216 319
rect 171 314 176 317
rect 104 310 118 314
rect 84 308 87 310
rect 89 308 91 310
rect 84 306 91 308
rect 109 309 118 310
rect 109 307 111 309
rect 113 307 118 309
rect 36 302 38 304
rect 40 302 42 304
rect 36 300 42 302
rect 66 300 73 306
rect 109 305 118 307
rect 120 312 128 314
rect 120 310 123 312
rect 125 310 128 312
rect 120 305 128 310
rect 130 310 138 314
rect 130 308 133 310
rect 135 308 138 310
rect 130 305 138 308
rect 66 298 68 300
rect 70 298 73 300
rect 66 296 73 298
rect 133 302 138 305
rect 140 302 145 314
rect 147 302 155 314
rect 169 312 176 314
rect 169 310 171 312
rect 173 310 176 312
rect 169 308 176 310
rect 178 308 189 317
rect 180 306 189 308
rect 191 306 196 317
rect 198 312 203 317
rect 209 315 211 317
rect 213 315 216 317
rect 209 313 216 315
rect 198 310 205 312
rect 211 310 216 313
rect 218 314 223 319
rect 218 310 232 314
rect 198 308 201 310
rect 203 308 205 310
rect 198 306 205 308
rect 223 309 232 310
rect 223 307 225 309
rect 227 307 232 309
rect 149 300 155 302
rect 149 298 151 300
rect 153 298 155 300
rect 149 296 155 298
rect 180 300 187 306
rect 223 305 232 307
rect 234 312 242 314
rect 234 310 237 312
rect 239 310 242 312
rect 234 305 242 310
rect 244 310 252 314
rect 244 308 247 310
rect 249 308 252 310
rect 244 305 252 308
rect 180 298 182 300
rect 184 298 187 300
rect 180 296 187 298
rect 247 302 252 305
rect 254 302 259 314
rect 261 302 269 314
rect 282 312 287 317
rect 280 310 287 312
rect 280 308 282 310
rect 284 308 287 310
rect 280 306 287 308
rect 289 306 294 317
rect 296 308 307 317
rect 309 314 314 317
rect 309 312 316 314
rect 368 313 373 314
rect 309 310 312 312
rect 314 310 316 312
rect 309 308 316 310
rect 322 311 329 313
rect 322 309 324 311
rect 326 309 329 311
rect 296 306 305 308
rect 263 300 269 302
rect 263 298 265 300
rect 267 298 269 300
rect 263 296 269 298
rect 298 300 305 306
rect 322 307 329 309
rect 331 311 339 313
rect 331 309 334 311
rect 336 309 339 311
rect 331 307 339 309
rect 298 298 301 300
rect 303 298 305 300
rect 298 296 305 298
rect 333 305 339 307
rect 341 305 346 313
rect 348 309 356 313
rect 348 307 351 309
rect 353 307 356 309
rect 348 305 356 307
rect 358 305 363 313
rect 365 309 373 313
rect 365 307 368 309
rect 370 307 373 309
rect 365 305 373 307
rect 375 312 382 314
rect 375 310 378 312
rect 380 310 382 312
rect 375 308 382 310
rect 389 312 396 314
rect 389 310 391 312
rect 393 310 396 312
rect 389 308 396 310
rect 375 305 380 308
rect 391 305 396 308
rect 398 313 403 314
rect 398 309 406 313
rect 398 307 401 309
rect 403 307 406 309
rect 398 305 406 307
rect 408 305 413 313
rect 415 309 423 313
rect 415 307 418 309
rect 420 307 423 309
rect 415 305 423 307
rect 425 305 430 313
rect 432 311 440 313
rect 432 309 435 311
rect 437 309 440 311
rect 432 307 440 309
rect 442 311 449 313
rect 442 309 445 311
rect 447 309 449 311
rect 442 307 449 309
rect 456 312 463 314
rect 456 310 458 312
rect 460 310 463 312
rect 456 308 463 310
rect 432 305 438 307
rect 458 305 463 308
rect 465 313 470 314
rect 522 317 529 319
rect 522 315 524 317
rect 526 315 529 317
rect 522 313 529 315
rect 465 309 473 313
rect 465 307 468 309
rect 470 307 473 309
rect 465 305 473 307
rect 475 305 480 313
rect 482 309 490 313
rect 482 307 485 309
rect 487 307 490 309
rect 482 305 490 307
rect 492 305 497 313
rect 499 311 507 313
rect 499 309 502 311
rect 504 309 507 311
rect 499 307 507 309
rect 509 311 516 313
rect 509 309 512 311
rect 514 309 516 311
rect 524 310 529 313
rect 531 313 539 319
rect 541 317 549 319
rect 541 315 544 317
rect 546 315 549 317
rect 541 313 549 315
rect 551 313 558 319
rect 610 314 615 319
rect 531 310 537 313
rect 509 307 516 309
rect 499 305 505 307
rect 533 306 537 310
rect 553 306 558 313
rect 533 304 539 306
rect 533 302 535 304
rect 537 302 539 304
rect 533 300 539 302
rect 552 304 558 306
rect 552 302 554 304
rect 556 302 558 304
rect 552 300 558 302
rect 564 302 572 314
rect 574 302 579 314
rect 581 310 589 314
rect 581 308 584 310
rect 586 308 589 310
rect 581 305 589 308
rect 591 312 599 314
rect 591 310 594 312
rect 596 310 599 312
rect 591 305 599 310
rect 601 310 615 314
rect 617 317 624 319
rect 617 315 620 317
rect 622 315 624 317
rect 617 313 624 315
rect 617 310 622 313
rect 601 309 610 310
rect 601 307 606 309
rect 608 307 610 309
rect 601 305 610 307
rect 581 302 586 305
rect 564 300 570 302
rect 564 298 566 300
rect 568 298 570 300
rect 564 296 570 298
rect 17 284 23 286
rect 17 282 19 284
rect 21 282 23 284
rect 17 280 23 282
rect 36 284 42 286
rect 66 288 73 290
rect 66 286 68 288
rect 70 286 73 288
rect 36 282 38 284
rect 40 282 42 284
rect 36 280 42 282
rect 17 276 21 280
rect 8 273 13 276
rect 6 271 13 273
rect 6 269 8 271
rect 10 269 13 271
rect 6 267 13 269
rect 15 273 21 276
rect 37 273 42 280
rect 66 280 73 286
rect 149 288 155 290
rect 149 286 151 288
rect 153 286 155 288
rect 149 284 155 286
rect 180 288 187 290
rect 180 286 182 288
rect 184 286 187 288
rect 133 281 138 284
rect 66 278 75 280
rect 15 267 23 273
rect 25 271 33 273
rect 25 269 28 271
rect 30 269 33 271
rect 25 267 33 269
rect 35 267 42 273
rect 55 276 62 278
rect 55 274 57 276
rect 59 274 62 276
rect 55 272 62 274
rect 57 269 62 272
rect 64 269 75 278
rect 77 269 82 280
rect 84 278 91 280
rect 84 276 87 278
rect 89 276 91 278
rect 109 279 118 281
rect 109 277 111 279
rect 113 277 118 279
rect 109 276 118 277
rect 84 274 91 276
rect 84 269 89 274
rect 97 273 102 276
rect 95 271 102 273
rect 95 269 97 271
rect 99 269 102 271
rect 95 267 102 269
rect 104 272 118 276
rect 120 276 128 281
rect 120 274 123 276
rect 125 274 128 276
rect 120 272 128 274
rect 130 278 138 281
rect 130 276 133 278
rect 135 276 138 278
rect 130 272 138 276
rect 140 272 145 284
rect 147 272 155 284
rect 180 280 187 286
rect 263 288 269 290
rect 263 286 265 288
rect 267 286 269 288
rect 263 284 269 286
rect 298 288 305 290
rect 298 286 301 288
rect 303 286 305 288
rect 247 281 252 284
rect 180 278 189 280
rect 169 276 176 278
rect 169 274 171 276
rect 173 274 176 276
rect 169 272 176 274
rect 104 267 109 272
rect 171 269 176 272
rect 178 269 189 278
rect 191 269 196 280
rect 198 278 205 280
rect 198 276 201 278
rect 203 276 205 278
rect 223 279 232 281
rect 223 277 225 279
rect 227 277 232 279
rect 223 276 232 277
rect 198 274 205 276
rect 198 269 203 274
rect 211 273 216 276
rect 209 271 216 273
rect 209 269 211 271
rect 213 269 216 271
rect 209 267 216 269
rect 218 272 232 276
rect 234 276 242 281
rect 234 274 237 276
rect 239 274 242 276
rect 234 272 242 274
rect 244 278 252 281
rect 244 276 247 278
rect 249 276 252 278
rect 244 272 252 276
rect 254 272 259 284
rect 261 272 269 284
rect 298 280 305 286
rect 280 278 287 280
rect 280 276 282 278
rect 284 276 287 278
rect 280 274 287 276
rect 218 267 223 272
rect 282 269 287 274
rect 289 269 294 280
rect 296 278 305 280
rect 333 279 339 281
rect 296 269 307 278
rect 309 276 316 278
rect 309 274 312 276
rect 314 274 316 276
rect 309 272 316 274
rect 322 277 329 279
rect 322 275 324 277
rect 326 275 329 277
rect 322 273 329 275
rect 331 277 339 279
rect 331 275 334 277
rect 336 275 339 277
rect 331 273 339 275
rect 341 273 346 281
rect 348 279 356 281
rect 348 277 351 279
rect 353 277 356 279
rect 348 273 356 277
rect 358 273 363 281
rect 365 279 373 281
rect 365 277 368 279
rect 370 277 373 279
rect 365 273 373 277
rect 309 269 314 272
rect 368 272 373 273
rect 375 278 380 281
rect 391 278 396 281
rect 375 276 382 278
rect 375 274 378 276
rect 380 274 382 276
rect 375 272 382 274
rect 389 276 396 278
rect 389 274 391 276
rect 393 274 396 276
rect 389 272 396 274
rect 398 279 406 281
rect 398 277 401 279
rect 403 277 406 279
rect 398 273 406 277
rect 408 273 413 281
rect 415 279 423 281
rect 415 277 418 279
rect 420 277 423 279
rect 415 273 423 277
rect 425 273 430 281
rect 432 279 438 281
rect 432 277 440 279
rect 432 275 435 277
rect 437 275 440 277
rect 432 273 440 275
rect 442 277 449 279
rect 458 278 463 281
rect 442 275 445 277
rect 447 275 449 277
rect 442 273 449 275
rect 456 276 463 278
rect 456 274 458 276
rect 460 274 463 276
rect 398 272 403 273
rect 456 272 463 274
rect 465 279 473 281
rect 465 277 468 279
rect 470 277 473 279
rect 465 273 473 277
rect 475 273 480 281
rect 482 279 490 281
rect 482 277 485 279
rect 487 277 490 279
rect 482 273 490 277
rect 492 273 497 281
rect 499 279 505 281
rect 564 288 570 290
rect 564 286 566 288
rect 568 286 570 288
rect 533 284 539 286
rect 533 282 535 284
rect 537 282 539 284
rect 499 277 507 279
rect 499 275 502 277
rect 504 275 507 277
rect 499 273 507 275
rect 509 277 516 279
rect 509 275 512 277
rect 514 275 516 277
rect 533 280 539 282
rect 552 284 558 286
rect 552 282 554 284
rect 556 282 558 284
rect 552 280 558 282
rect 533 276 537 280
rect 509 273 516 275
rect 524 273 529 276
rect 465 272 470 273
rect 522 271 529 273
rect 522 269 524 271
rect 526 269 529 271
rect 522 267 529 269
rect 531 273 537 276
rect 553 273 558 280
rect 531 267 539 273
rect 541 271 549 273
rect 541 269 544 271
rect 546 269 549 271
rect 541 267 549 269
rect 551 267 558 273
rect 564 284 570 286
rect 564 272 572 284
rect 574 272 579 284
rect 581 281 586 284
rect 581 278 589 281
rect 581 276 584 278
rect 586 276 589 278
rect 581 272 589 276
rect 591 276 599 281
rect 591 274 594 276
rect 596 274 599 276
rect 591 272 599 274
rect 601 279 610 281
rect 601 277 606 279
rect 608 277 610 279
rect 601 276 610 277
rect 601 272 615 276
rect 610 267 615 272
rect 617 273 622 276
rect 617 271 624 273
rect 617 269 620 271
rect 622 269 624 271
rect 617 267 624 269
rect 6 173 13 175
rect 6 171 8 173
rect 10 171 13 173
rect 6 169 13 171
rect 8 166 13 169
rect 15 169 23 175
rect 25 173 33 175
rect 25 171 28 173
rect 30 171 33 173
rect 25 169 33 171
rect 35 169 42 175
rect 95 173 102 175
rect 57 170 62 173
rect 15 166 21 169
rect 17 162 21 166
rect 37 162 42 169
rect 55 168 62 170
rect 55 166 57 168
rect 59 166 62 168
rect 55 164 62 166
rect 64 164 75 173
rect 17 160 23 162
rect 17 158 19 160
rect 21 158 23 160
rect 17 156 23 158
rect 36 160 42 162
rect 66 162 75 164
rect 77 162 82 173
rect 84 168 89 173
rect 95 171 97 173
rect 99 171 102 173
rect 95 169 102 171
rect 84 166 91 168
rect 97 166 102 169
rect 104 170 109 175
rect 209 173 216 175
rect 171 170 176 173
rect 104 166 118 170
rect 84 164 87 166
rect 89 164 91 166
rect 84 162 91 164
rect 109 165 118 166
rect 109 163 111 165
rect 113 163 118 165
rect 36 158 38 160
rect 40 158 42 160
rect 36 156 42 158
rect 66 156 73 162
rect 109 161 118 163
rect 120 168 128 170
rect 120 166 123 168
rect 125 166 128 168
rect 120 161 128 166
rect 130 166 138 170
rect 130 164 133 166
rect 135 164 138 166
rect 130 161 138 164
rect 66 154 68 156
rect 70 154 73 156
rect 66 152 73 154
rect 133 158 138 161
rect 140 158 145 170
rect 147 158 155 170
rect 169 168 176 170
rect 169 166 171 168
rect 173 166 176 168
rect 169 164 176 166
rect 178 164 189 173
rect 180 162 189 164
rect 191 162 196 173
rect 198 168 203 173
rect 209 171 211 173
rect 213 171 216 173
rect 209 169 216 171
rect 198 166 205 168
rect 211 166 216 169
rect 218 170 223 175
rect 218 166 232 170
rect 198 164 201 166
rect 203 164 205 166
rect 198 162 205 164
rect 223 165 232 166
rect 223 163 225 165
rect 227 163 232 165
rect 149 156 155 158
rect 149 154 151 156
rect 153 154 155 156
rect 149 152 155 154
rect 180 156 187 162
rect 223 161 232 163
rect 234 168 242 170
rect 234 166 237 168
rect 239 166 242 168
rect 234 161 242 166
rect 244 166 252 170
rect 244 164 247 166
rect 249 164 252 166
rect 244 161 252 164
rect 180 154 182 156
rect 184 154 187 156
rect 180 152 187 154
rect 247 158 252 161
rect 254 158 259 170
rect 261 158 269 170
rect 282 168 287 173
rect 280 166 287 168
rect 280 164 282 166
rect 284 164 287 166
rect 280 162 287 164
rect 289 162 294 173
rect 296 164 307 173
rect 309 170 314 173
rect 309 168 316 170
rect 368 169 373 170
rect 309 166 312 168
rect 314 166 316 168
rect 309 164 316 166
rect 322 167 329 169
rect 322 165 324 167
rect 326 165 329 167
rect 296 162 305 164
rect 263 156 269 158
rect 263 154 265 156
rect 267 154 269 156
rect 263 152 269 154
rect 298 156 305 162
rect 322 163 329 165
rect 331 167 339 169
rect 331 165 334 167
rect 336 165 339 167
rect 331 163 339 165
rect 298 154 301 156
rect 303 154 305 156
rect 298 152 305 154
rect 333 161 339 163
rect 341 161 346 169
rect 348 165 356 169
rect 348 163 351 165
rect 353 163 356 165
rect 348 161 356 163
rect 358 161 363 169
rect 365 165 373 169
rect 365 163 368 165
rect 370 163 373 165
rect 365 161 373 163
rect 375 168 382 170
rect 375 166 378 168
rect 380 166 382 168
rect 375 164 382 166
rect 389 168 396 170
rect 389 166 391 168
rect 393 166 396 168
rect 389 164 396 166
rect 375 161 380 164
rect 391 161 396 164
rect 398 169 403 170
rect 398 165 406 169
rect 398 163 401 165
rect 403 163 406 165
rect 398 161 406 163
rect 408 161 413 169
rect 415 165 423 169
rect 415 163 418 165
rect 420 163 423 165
rect 415 161 423 163
rect 425 161 430 169
rect 432 167 440 169
rect 432 165 435 167
rect 437 165 440 167
rect 432 163 440 165
rect 442 167 449 169
rect 442 165 445 167
rect 447 165 449 167
rect 442 163 449 165
rect 456 168 463 170
rect 456 166 458 168
rect 460 166 463 168
rect 456 164 463 166
rect 432 161 438 163
rect 458 161 463 164
rect 465 169 470 170
rect 522 173 529 175
rect 522 171 524 173
rect 526 171 529 173
rect 522 169 529 171
rect 465 165 473 169
rect 465 163 468 165
rect 470 163 473 165
rect 465 161 473 163
rect 475 161 480 169
rect 482 165 490 169
rect 482 163 485 165
rect 487 163 490 165
rect 482 161 490 163
rect 492 161 497 169
rect 499 167 507 169
rect 499 165 502 167
rect 504 165 507 167
rect 499 163 507 165
rect 509 167 516 169
rect 509 165 512 167
rect 514 165 516 167
rect 524 166 529 169
rect 531 169 539 175
rect 541 173 549 175
rect 541 171 544 173
rect 546 171 549 173
rect 541 169 549 171
rect 551 169 558 175
rect 610 170 615 175
rect 531 166 537 169
rect 509 163 516 165
rect 499 161 505 163
rect 533 162 537 166
rect 553 162 558 169
rect 533 160 539 162
rect 533 158 535 160
rect 537 158 539 160
rect 533 156 539 158
rect 552 160 558 162
rect 552 158 554 160
rect 556 158 558 160
rect 552 156 558 158
rect 564 158 572 170
rect 574 158 579 170
rect 581 166 589 170
rect 581 164 584 166
rect 586 164 589 166
rect 581 161 589 164
rect 591 168 599 170
rect 591 166 594 168
rect 596 166 599 168
rect 591 161 599 166
rect 601 166 615 170
rect 617 173 624 175
rect 617 171 620 173
rect 622 171 624 173
rect 617 169 624 171
rect 617 166 622 169
rect 601 165 610 166
rect 601 163 606 165
rect 608 163 610 165
rect 601 161 610 163
rect 581 158 586 161
rect 564 156 570 158
rect 564 154 566 156
rect 568 154 570 156
rect 564 152 570 154
rect 17 140 23 142
rect 17 138 19 140
rect 21 138 23 140
rect 17 136 23 138
rect 36 140 42 142
rect 66 144 73 146
rect 66 142 68 144
rect 70 142 73 144
rect 36 138 38 140
rect 40 138 42 140
rect 36 136 42 138
rect 17 132 21 136
rect 8 129 13 132
rect 6 127 13 129
rect 6 125 8 127
rect 10 125 13 127
rect 6 123 13 125
rect 15 129 21 132
rect 37 129 42 136
rect 66 136 73 142
rect 149 144 155 146
rect 149 142 151 144
rect 153 142 155 144
rect 149 140 155 142
rect 180 144 187 146
rect 180 142 182 144
rect 184 142 187 144
rect 133 137 138 140
rect 66 134 75 136
rect 15 123 23 129
rect 25 127 33 129
rect 25 125 28 127
rect 30 125 33 127
rect 25 123 33 125
rect 35 123 42 129
rect 55 132 62 134
rect 55 130 57 132
rect 59 130 62 132
rect 55 128 62 130
rect 57 125 62 128
rect 64 125 75 134
rect 77 125 82 136
rect 84 134 91 136
rect 84 132 87 134
rect 89 132 91 134
rect 109 135 118 137
rect 109 133 111 135
rect 113 133 118 135
rect 109 132 118 133
rect 84 130 91 132
rect 84 125 89 130
rect 97 129 102 132
rect 95 127 102 129
rect 95 125 97 127
rect 99 125 102 127
rect 95 123 102 125
rect 104 128 118 132
rect 120 132 128 137
rect 120 130 123 132
rect 125 130 128 132
rect 120 128 128 130
rect 130 134 138 137
rect 130 132 133 134
rect 135 132 138 134
rect 130 128 138 132
rect 140 128 145 140
rect 147 128 155 140
rect 180 136 187 142
rect 263 144 269 146
rect 263 142 265 144
rect 267 142 269 144
rect 263 140 269 142
rect 298 144 305 146
rect 298 142 301 144
rect 303 142 305 144
rect 247 137 252 140
rect 180 134 189 136
rect 169 132 176 134
rect 169 130 171 132
rect 173 130 176 132
rect 169 128 176 130
rect 104 123 109 128
rect 171 125 176 128
rect 178 125 189 134
rect 191 125 196 136
rect 198 134 205 136
rect 198 132 201 134
rect 203 132 205 134
rect 223 135 232 137
rect 223 133 225 135
rect 227 133 232 135
rect 223 132 232 133
rect 198 130 205 132
rect 198 125 203 130
rect 211 129 216 132
rect 209 127 216 129
rect 209 125 211 127
rect 213 125 216 127
rect 209 123 216 125
rect 218 128 232 132
rect 234 132 242 137
rect 234 130 237 132
rect 239 130 242 132
rect 234 128 242 130
rect 244 134 252 137
rect 244 132 247 134
rect 249 132 252 134
rect 244 128 252 132
rect 254 128 259 140
rect 261 128 269 140
rect 298 136 305 142
rect 280 134 287 136
rect 280 132 282 134
rect 284 132 287 134
rect 280 130 287 132
rect 218 123 223 128
rect 282 125 287 130
rect 289 125 294 136
rect 296 134 305 136
rect 333 135 339 137
rect 296 125 307 134
rect 309 132 316 134
rect 309 130 312 132
rect 314 130 316 132
rect 309 128 316 130
rect 322 133 329 135
rect 322 131 324 133
rect 326 131 329 133
rect 322 129 329 131
rect 331 133 339 135
rect 331 131 334 133
rect 336 131 339 133
rect 331 129 339 131
rect 341 129 346 137
rect 348 135 356 137
rect 348 133 351 135
rect 353 133 356 135
rect 348 129 356 133
rect 358 129 363 137
rect 365 135 373 137
rect 365 133 368 135
rect 370 133 373 135
rect 365 129 373 133
rect 309 125 314 128
rect 368 128 373 129
rect 375 134 380 137
rect 391 134 396 137
rect 375 132 382 134
rect 375 130 378 132
rect 380 130 382 132
rect 375 128 382 130
rect 389 132 396 134
rect 389 130 391 132
rect 393 130 396 132
rect 389 128 396 130
rect 398 135 406 137
rect 398 133 401 135
rect 403 133 406 135
rect 398 129 406 133
rect 408 129 413 137
rect 415 135 423 137
rect 415 133 418 135
rect 420 133 423 135
rect 415 129 423 133
rect 425 129 430 137
rect 432 135 438 137
rect 432 133 440 135
rect 432 131 435 133
rect 437 131 440 133
rect 432 129 440 131
rect 442 133 449 135
rect 458 134 463 137
rect 442 131 445 133
rect 447 131 449 133
rect 442 129 449 131
rect 456 132 463 134
rect 456 130 458 132
rect 460 130 463 132
rect 398 128 403 129
rect 456 128 463 130
rect 465 135 473 137
rect 465 133 468 135
rect 470 133 473 135
rect 465 129 473 133
rect 475 129 480 137
rect 482 135 490 137
rect 482 133 485 135
rect 487 133 490 135
rect 482 129 490 133
rect 492 129 497 137
rect 499 135 505 137
rect 564 144 570 146
rect 564 142 566 144
rect 568 142 570 144
rect 533 140 539 142
rect 533 138 535 140
rect 537 138 539 140
rect 499 133 507 135
rect 499 131 502 133
rect 504 131 507 133
rect 499 129 507 131
rect 509 133 516 135
rect 509 131 512 133
rect 514 131 516 133
rect 533 136 539 138
rect 552 140 558 142
rect 552 138 554 140
rect 556 138 558 140
rect 552 136 558 138
rect 533 132 537 136
rect 509 129 516 131
rect 524 129 529 132
rect 465 128 470 129
rect 522 127 529 129
rect 522 125 524 127
rect 526 125 529 127
rect 522 123 529 125
rect 531 129 537 132
rect 553 129 558 136
rect 531 123 539 129
rect 541 127 549 129
rect 541 125 544 127
rect 546 125 549 127
rect 541 123 549 125
rect 551 123 558 129
rect 564 140 570 142
rect 564 128 572 140
rect 574 128 579 140
rect 581 137 586 140
rect 581 134 589 137
rect 581 132 584 134
rect 586 132 589 134
rect 581 128 589 132
rect 591 132 599 137
rect 591 130 594 132
rect 596 130 599 132
rect 591 128 599 130
rect 601 135 610 137
rect 601 133 606 135
rect 608 133 610 135
rect 601 132 610 133
rect 601 128 615 132
rect 610 123 615 128
rect 617 129 622 132
rect 617 127 624 129
rect 617 125 620 127
rect 622 125 624 127
rect 617 123 624 125
rect 6 29 13 31
rect 6 27 8 29
rect 10 27 13 29
rect 6 25 13 27
rect 8 22 13 25
rect 15 25 23 31
rect 25 29 33 31
rect 25 27 28 29
rect 30 27 33 29
rect 25 25 33 27
rect 35 25 42 31
rect 95 29 102 31
rect 57 26 62 29
rect 15 22 21 25
rect 17 18 21 22
rect 37 18 42 25
rect 55 24 62 26
rect 55 22 57 24
rect 59 22 62 24
rect 55 20 62 22
rect 64 20 75 29
rect 17 16 23 18
rect 17 14 19 16
rect 21 14 23 16
rect 17 12 23 14
rect 36 16 42 18
rect 66 18 75 20
rect 77 18 82 29
rect 84 24 89 29
rect 95 27 97 29
rect 99 27 102 29
rect 95 25 102 27
rect 84 22 91 24
rect 97 22 102 25
rect 104 26 109 31
rect 209 29 216 31
rect 171 26 176 29
rect 104 22 118 26
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 109 21 118 22
rect 109 19 111 21
rect 113 19 118 21
rect 36 14 38 16
rect 40 14 42 16
rect 36 12 42 14
rect 66 12 73 18
rect 109 17 118 19
rect 120 24 128 26
rect 120 22 123 24
rect 125 22 128 24
rect 120 17 128 22
rect 130 22 138 26
rect 130 20 133 22
rect 135 20 138 22
rect 130 17 138 20
rect 66 10 68 12
rect 70 10 73 12
rect 66 8 73 10
rect 133 14 138 17
rect 140 14 145 26
rect 147 14 155 26
rect 169 24 176 26
rect 169 22 171 24
rect 173 22 176 24
rect 169 20 176 22
rect 178 20 189 29
rect 180 18 189 20
rect 191 18 196 29
rect 198 24 203 29
rect 209 27 211 29
rect 213 27 216 29
rect 209 25 216 27
rect 198 22 205 24
rect 211 22 216 25
rect 218 26 223 31
rect 218 22 232 26
rect 198 20 201 22
rect 203 20 205 22
rect 198 18 205 20
rect 223 21 232 22
rect 223 19 225 21
rect 227 19 232 21
rect 149 12 155 14
rect 149 10 151 12
rect 153 10 155 12
rect 149 8 155 10
rect 180 12 187 18
rect 223 17 232 19
rect 234 24 242 26
rect 234 22 237 24
rect 239 22 242 24
rect 234 17 242 22
rect 244 22 252 26
rect 244 20 247 22
rect 249 20 252 22
rect 244 17 252 20
rect 180 10 182 12
rect 184 10 187 12
rect 180 8 187 10
rect 247 14 252 17
rect 254 14 259 26
rect 261 14 269 26
rect 282 24 287 29
rect 280 22 287 24
rect 280 20 282 22
rect 284 20 287 22
rect 280 18 287 20
rect 289 18 294 29
rect 296 20 307 29
rect 309 26 314 29
rect 309 24 316 26
rect 368 25 373 26
rect 309 22 312 24
rect 314 22 316 24
rect 309 20 316 22
rect 322 23 329 25
rect 322 21 324 23
rect 326 21 329 23
rect 296 18 305 20
rect 263 12 269 14
rect 263 10 265 12
rect 267 10 269 12
rect 263 8 269 10
rect 298 12 305 18
rect 322 19 329 21
rect 331 23 339 25
rect 331 21 334 23
rect 336 21 339 23
rect 331 19 339 21
rect 298 10 301 12
rect 303 10 305 12
rect 298 8 305 10
rect 333 17 339 19
rect 341 17 346 25
rect 348 21 356 25
rect 348 19 351 21
rect 353 19 356 21
rect 348 17 356 19
rect 358 17 363 25
rect 365 21 373 25
rect 365 19 368 21
rect 370 19 373 21
rect 365 17 373 19
rect 375 24 382 26
rect 375 22 378 24
rect 380 22 382 24
rect 375 20 382 22
rect 389 24 396 26
rect 389 22 391 24
rect 393 22 396 24
rect 389 20 396 22
rect 375 17 380 20
rect 391 17 396 20
rect 398 25 403 26
rect 398 21 406 25
rect 398 19 401 21
rect 403 19 406 21
rect 398 17 406 19
rect 408 17 413 25
rect 415 21 423 25
rect 415 19 418 21
rect 420 19 423 21
rect 415 17 423 19
rect 425 17 430 25
rect 432 23 440 25
rect 432 21 435 23
rect 437 21 440 23
rect 432 19 440 21
rect 442 23 449 25
rect 442 21 445 23
rect 447 21 449 23
rect 442 19 449 21
rect 456 24 463 26
rect 456 22 458 24
rect 460 22 463 24
rect 456 20 463 22
rect 432 17 438 19
rect 458 17 463 20
rect 465 25 470 26
rect 522 29 529 31
rect 522 27 524 29
rect 526 27 529 29
rect 522 25 529 27
rect 465 21 473 25
rect 465 19 468 21
rect 470 19 473 21
rect 465 17 473 19
rect 475 17 480 25
rect 482 21 490 25
rect 482 19 485 21
rect 487 19 490 21
rect 482 17 490 19
rect 492 17 497 25
rect 499 23 507 25
rect 499 21 502 23
rect 504 21 507 23
rect 499 19 507 21
rect 509 23 516 25
rect 509 21 512 23
rect 514 21 516 23
rect 524 22 529 25
rect 531 25 539 31
rect 541 29 549 31
rect 541 27 544 29
rect 546 27 549 29
rect 541 25 549 27
rect 551 25 558 31
rect 610 26 615 31
rect 531 22 537 25
rect 509 19 516 21
rect 499 17 505 19
rect 533 18 537 22
rect 553 18 558 25
rect 533 16 539 18
rect 533 14 535 16
rect 537 14 539 16
rect 533 12 539 14
rect 552 16 558 18
rect 552 14 554 16
rect 556 14 558 16
rect 552 12 558 14
rect 564 14 572 26
rect 574 14 579 26
rect 581 22 589 26
rect 581 20 584 22
rect 586 20 589 22
rect 581 17 589 20
rect 591 24 599 26
rect 591 22 594 24
rect 596 22 599 24
rect 591 17 599 22
rect 601 22 615 26
rect 617 29 624 31
rect 617 27 620 29
rect 622 27 624 29
rect 617 25 624 27
rect 617 22 622 25
rect 601 21 610 22
rect 601 19 606 21
rect 608 19 610 21
rect 601 17 610 19
rect 581 14 586 17
rect 564 12 570 14
rect 564 10 566 12
rect 568 10 570 12
rect 564 8 570 10
<< pdif >>
rect 8 538 13 543
rect 6 536 13 538
rect 6 534 8 536
rect 10 534 13 536
rect 6 529 13 534
rect 6 527 8 529
rect 10 527 13 529
rect 6 525 13 527
rect 15 536 23 543
rect 55 540 62 542
rect 55 538 57 540
rect 59 538 62 540
rect 15 525 26 536
rect 17 519 26 525
rect 17 517 19 519
rect 21 517 26 519
rect 17 515 26 517
rect 28 515 33 536
rect 35 528 40 536
rect 55 533 62 538
rect 55 531 57 533
rect 59 531 62 533
rect 55 529 62 531
rect 35 526 42 528
rect 35 524 38 526
rect 40 524 42 526
rect 57 524 62 529
rect 64 535 70 542
rect 103 540 110 542
rect 103 538 105 540
rect 107 538 110 540
rect 103 536 110 538
rect 64 528 72 535
rect 64 526 67 528
rect 69 526 72 528
rect 64 524 72 526
rect 35 522 42 524
rect 35 515 40 522
rect 66 522 72 524
rect 74 533 82 535
rect 74 531 77 533
rect 79 531 82 533
rect 74 526 82 531
rect 74 524 77 526
rect 79 524 82 526
rect 74 522 82 524
rect 84 526 91 535
rect 84 524 87 526
rect 89 524 91 526
rect 84 522 91 524
rect 105 515 110 536
rect 112 526 126 542
rect 112 524 115 526
rect 117 524 126 526
rect 128 540 136 542
rect 128 538 131 540
rect 133 538 136 540
rect 128 533 136 538
rect 128 531 131 533
rect 133 531 136 533
rect 128 524 136 531
rect 138 533 146 542
rect 138 531 141 533
rect 143 531 146 533
rect 138 524 146 531
rect 112 519 124 524
rect 112 517 115 519
rect 117 517 124 519
rect 112 515 124 517
rect 141 515 146 524
rect 148 527 153 542
rect 169 540 176 542
rect 169 538 171 540
rect 173 538 176 540
rect 169 533 176 538
rect 169 531 171 533
rect 173 531 176 533
rect 169 529 176 531
rect 148 525 155 527
rect 148 523 151 525
rect 153 523 155 525
rect 171 524 176 529
rect 178 535 184 542
rect 217 540 224 542
rect 217 538 219 540
rect 221 538 224 540
rect 217 536 224 538
rect 178 528 186 535
rect 178 526 181 528
rect 183 526 186 528
rect 178 524 186 526
rect 148 521 155 523
rect 148 515 153 521
rect 180 522 186 524
rect 188 533 196 535
rect 188 531 191 533
rect 193 531 196 533
rect 188 526 196 531
rect 188 524 191 526
rect 193 524 196 526
rect 188 522 196 524
rect 198 526 205 535
rect 198 524 201 526
rect 203 524 205 526
rect 198 522 205 524
rect 219 515 224 536
rect 226 526 240 542
rect 226 524 229 526
rect 231 524 240 526
rect 242 540 250 542
rect 242 538 245 540
rect 247 538 250 540
rect 242 533 250 538
rect 242 531 245 533
rect 247 531 250 533
rect 242 524 250 531
rect 252 533 260 542
rect 252 531 255 533
rect 257 531 260 533
rect 252 524 260 531
rect 226 519 238 524
rect 226 517 229 519
rect 231 517 238 519
rect 226 515 238 517
rect 255 515 260 524
rect 262 527 267 542
rect 301 535 307 542
rect 262 525 269 527
rect 262 523 265 525
rect 267 523 269 525
rect 262 521 269 523
rect 280 526 287 535
rect 280 524 282 526
rect 284 524 287 526
rect 280 522 287 524
rect 289 533 297 535
rect 289 531 292 533
rect 294 531 297 533
rect 289 526 297 531
rect 289 524 292 526
rect 294 524 297 526
rect 289 522 297 524
rect 299 528 307 535
rect 299 526 302 528
rect 304 526 307 528
rect 299 524 307 526
rect 309 540 316 542
rect 309 538 312 540
rect 314 538 316 540
rect 309 533 316 538
rect 322 541 329 543
rect 322 539 324 541
rect 326 539 329 541
rect 322 537 329 539
rect 324 535 329 537
rect 331 535 337 543
rect 309 531 312 533
rect 314 531 316 533
rect 309 529 316 531
rect 333 531 337 535
rect 368 531 373 533
rect 309 524 314 529
rect 333 527 339 531
rect 299 522 305 524
rect 262 515 267 521
rect 332 519 339 527
rect 332 517 334 519
rect 336 517 339 519
rect 332 515 339 517
rect 341 515 346 531
rect 348 529 356 531
rect 348 527 351 529
rect 353 527 356 529
rect 348 515 356 527
rect 358 515 363 531
rect 365 519 373 531
rect 365 517 368 519
rect 370 517 373 519
rect 365 515 373 517
rect 375 528 380 533
rect 391 528 396 533
rect 375 526 382 528
rect 375 524 378 526
rect 380 524 382 526
rect 375 522 382 524
rect 389 526 396 528
rect 389 524 391 526
rect 393 524 396 526
rect 389 522 396 524
rect 375 515 380 522
rect 391 515 396 522
rect 398 531 403 533
rect 434 535 440 543
rect 442 541 449 543
rect 442 539 445 541
rect 447 539 449 541
rect 442 537 449 539
rect 442 535 447 537
rect 434 531 438 535
rect 398 519 406 531
rect 398 517 401 519
rect 403 517 406 519
rect 398 515 406 517
rect 408 515 413 531
rect 415 529 423 531
rect 415 527 418 529
rect 420 527 423 529
rect 415 515 423 527
rect 425 515 430 531
rect 432 527 438 531
rect 458 528 463 533
rect 432 519 439 527
rect 456 526 463 528
rect 456 524 458 526
rect 460 524 463 526
rect 456 522 463 524
rect 432 517 435 519
rect 437 517 439 519
rect 432 515 439 517
rect 458 515 463 522
rect 465 531 470 533
rect 501 535 507 543
rect 509 541 516 543
rect 509 539 512 541
rect 514 539 516 541
rect 509 537 516 539
rect 524 538 529 543
rect 509 535 514 537
rect 522 536 529 538
rect 501 531 505 535
rect 465 519 473 531
rect 465 517 468 519
rect 470 517 473 519
rect 465 515 473 517
rect 475 515 480 531
rect 482 529 490 531
rect 482 527 485 529
rect 487 527 490 529
rect 482 515 490 527
rect 492 515 497 531
rect 499 527 505 531
rect 522 534 524 536
rect 526 534 529 536
rect 499 519 506 527
rect 522 529 529 534
rect 522 527 524 529
rect 526 527 529 529
rect 522 525 529 527
rect 531 536 539 543
rect 531 525 542 536
rect 499 517 502 519
rect 504 517 506 519
rect 533 519 542 525
rect 499 515 506 517
rect 533 517 535 519
rect 537 517 542 519
rect 533 515 542 517
rect 544 515 549 536
rect 551 528 556 536
rect 551 526 558 528
rect 566 527 571 542
rect 551 524 554 526
rect 556 524 558 526
rect 551 522 558 524
rect 564 525 571 527
rect 564 523 566 525
rect 568 523 571 525
rect 551 515 556 522
rect 564 521 571 523
rect 566 515 571 521
rect 573 533 581 542
rect 573 531 576 533
rect 578 531 581 533
rect 573 524 581 531
rect 583 540 591 542
rect 583 538 586 540
rect 588 538 591 540
rect 583 533 591 538
rect 583 531 586 533
rect 588 531 591 533
rect 583 524 591 531
rect 593 526 607 542
rect 593 524 602 526
rect 604 524 607 526
rect 573 515 578 524
rect 595 519 607 524
rect 595 517 602 519
rect 604 517 607 519
rect 595 515 607 517
rect 609 540 616 542
rect 609 538 612 540
rect 614 538 616 540
rect 609 536 616 538
rect 609 515 614 536
rect 17 501 26 503
rect 17 499 19 501
rect 21 499 26 501
rect 17 493 26 499
rect 6 491 13 493
rect 6 489 8 491
rect 10 489 13 491
rect 6 484 13 489
rect 6 482 8 484
rect 10 482 13 484
rect 6 480 13 482
rect 8 475 13 480
rect 15 482 26 493
rect 28 482 33 503
rect 35 496 40 503
rect 35 494 42 496
rect 66 494 72 496
rect 35 492 38 494
rect 40 492 42 494
rect 35 490 42 492
rect 35 482 40 490
rect 57 489 62 494
rect 55 487 62 489
rect 55 485 57 487
rect 59 485 62 487
rect 15 475 23 482
rect 55 480 62 485
rect 55 478 57 480
rect 59 478 62 480
rect 55 476 62 478
rect 64 492 72 494
rect 64 490 67 492
rect 69 490 72 492
rect 64 483 72 490
rect 74 494 82 496
rect 74 492 77 494
rect 79 492 82 494
rect 74 487 82 492
rect 74 485 77 487
rect 79 485 82 487
rect 74 483 82 485
rect 84 494 91 496
rect 84 492 87 494
rect 89 492 91 494
rect 84 483 91 492
rect 64 476 70 483
rect 105 482 110 503
rect 103 480 110 482
rect 103 478 105 480
rect 107 478 110 480
rect 103 476 110 478
rect 112 501 124 503
rect 112 499 115 501
rect 117 499 124 501
rect 112 494 124 499
rect 141 494 146 503
rect 112 492 115 494
rect 117 492 126 494
rect 112 476 126 492
rect 128 487 136 494
rect 128 485 131 487
rect 133 485 136 487
rect 128 480 136 485
rect 128 478 131 480
rect 133 478 136 480
rect 128 476 136 478
rect 138 487 146 494
rect 138 485 141 487
rect 143 485 146 487
rect 138 476 146 485
rect 148 497 153 503
rect 148 495 155 497
rect 148 493 151 495
rect 153 493 155 495
rect 180 494 186 496
rect 148 491 155 493
rect 148 476 153 491
rect 171 489 176 494
rect 169 487 176 489
rect 169 485 171 487
rect 173 485 176 487
rect 169 480 176 485
rect 169 478 171 480
rect 173 478 176 480
rect 169 476 176 478
rect 178 492 186 494
rect 178 490 181 492
rect 183 490 186 492
rect 178 483 186 490
rect 188 494 196 496
rect 188 492 191 494
rect 193 492 196 494
rect 188 487 196 492
rect 188 485 191 487
rect 193 485 196 487
rect 188 483 196 485
rect 198 494 205 496
rect 198 492 201 494
rect 203 492 205 494
rect 198 483 205 492
rect 178 476 184 483
rect 219 482 224 503
rect 217 480 224 482
rect 217 478 219 480
rect 221 478 224 480
rect 217 476 224 478
rect 226 501 238 503
rect 226 499 229 501
rect 231 499 238 501
rect 226 494 238 499
rect 255 494 260 503
rect 226 492 229 494
rect 231 492 240 494
rect 226 476 240 492
rect 242 487 250 494
rect 242 485 245 487
rect 247 485 250 487
rect 242 480 250 485
rect 242 478 245 480
rect 247 478 250 480
rect 242 476 250 478
rect 252 487 260 494
rect 252 485 255 487
rect 257 485 260 487
rect 252 476 260 485
rect 262 497 267 503
rect 262 495 269 497
rect 332 501 339 503
rect 332 499 334 501
rect 336 499 339 501
rect 262 493 265 495
rect 267 493 269 495
rect 262 491 269 493
rect 280 494 287 496
rect 280 492 282 494
rect 284 492 287 494
rect 262 476 267 491
rect 280 483 287 492
rect 289 494 297 496
rect 289 492 292 494
rect 294 492 297 494
rect 289 487 297 492
rect 289 485 292 487
rect 294 485 297 487
rect 289 483 297 485
rect 299 494 305 496
rect 299 492 307 494
rect 299 490 302 492
rect 304 490 307 492
rect 299 483 307 490
rect 301 476 307 483
rect 309 489 314 494
rect 332 491 339 499
rect 309 487 316 489
rect 309 485 312 487
rect 314 485 316 487
rect 309 480 316 485
rect 333 487 339 491
rect 341 487 346 503
rect 348 491 356 503
rect 348 489 351 491
rect 353 489 356 491
rect 348 487 356 489
rect 358 487 363 503
rect 365 501 373 503
rect 365 499 368 501
rect 370 499 373 501
rect 365 487 373 499
rect 333 483 337 487
rect 324 481 329 483
rect 309 478 312 480
rect 314 478 316 480
rect 309 476 316 478
rect 322 479 329 481
rect 322 477 324 479
rect 326 477 329 479
rect 322 475 329 477
rect 331 475 337 483
rect 368 485 373 487
rect 375 496 380 503
rect 391 496 396 503
rect 375 494 382 496
rect 375 492 378 494
rect 380 492 382 494
rect 375 490 382 492
rect 389 494 396 496
rect 389 492 391 494
rect 393 492 396 494
rect 389 490 396 492
rect 375 485 380 490
rect 391 485 396 490
rect 398 501 406 503
rect 398 499 401 501
rect 403 499 406 501
rect 398 487 406 499
rect 408 487 413 503
rect 415 491 423 503
rect 415 489 418 491
rect 420 489 423 491
rect 415 487 423 489
rect 425 487 430 503
rect 432 501 439 503
rect 432 499 435 501
rect 437 499 439 501
rect 432 491 439 499
rect 458 496 463 503
rect 456 494 463 496
rect 456 492 458 494
rect 460 492 463 494
rect 432 487 438 491
rect 456 490 463 492
rect 398 485 403 487
rect 434 483 438 487
rect 458 485 463 490
rect 465 501 473 503
rect 465 499 468 501
rect 470 499 473 501
rect 465 487 473 499
rect 475 487 480 503
rect 482 491 490 503
rect 482 489 485 491
rect 487 489 490 491
rect 482 487 490 489
rect 492 487 497 503
rect 499 501 506 503
rect 499 499 502 501
rect 504 499 506 501
rect 533 501 542 503
rect 499 491 506 499
rect 533 499 535 501
rect 537 499 542 501
rect 533 493 542 499
rect 499 487 505 491
rect 465 485 470 487
rect 434 475 440 483
rect 442 481 447 483
rect 442 479 449 481
rect 442 477 445 479
rect 447 477 449 479
rect 442 475 449 477
rect 501 483 505 487
rect 522 491 529 493
rect 522 489 524 491
rect 526 489 529 491
rect 522 484 529 489
rect 501 475 507 483
rect 509 481 514 483
rect 522 482 524 484
rect 526 482 529 484
rect 509 479 516 481
rect 522 480 529 482
rect 509 477 512 479
rect 514 477 516 479
rect 509 475 516 477
rect 524 475 529 480
rect 531 482 542 493
rect 544 482 549 503
rect 551 496 556 503
rect 566 497 571 503
rect 551 494 558 496
rect 551 492 554 494
rect 556 492 558 494
rect 551 490 558 492
rect 564 495 571 497
rect 564 493 566 495
rect 568 493 571 495
rect 564 491 571 493
rect 551 482 556 490
rect 531 475 539 482
rect 566 476 571 491
rect 573 494 578 503
rect 595 501 607 503
rect 595 499 602 501
rect 604 499 607 501
rect 595 494 607 499
rect 573 487 581 494
rect 573 485 576 487
rect 578 485 581 487
rect 573 476 581 485
rect 583 487 591 494
rect 583 485 586 487
rect 588 485 591 487
rect 583 480 591 485
rect 583 478 586 480
rect 588 478 591 480
rect 583 476 591 478
rect 593 492 602 494
rect 604 492 607 494
rect 593 476 607 492
rect 609 482 614 503
rect 609 480 616 482
rect 609 478 612 480
rect 614 478 616 480
rect 609 476 616 478
rect 8 394 13 399
rect 6 392 13 394
rect 6 390 8 392
rect 10 390 13 392
rect 6 385 13 390
rect 6 383 8 385
rect 10 383 13 385
rect 6 381 13 383
rect 15 392 23 399
rect 55 396 62 398
rect 55 394 57 396
rect 59 394 62 396
rect 15 381 26 392
rect 17 375 26 381
rect 17 373 19 375
rect 21 373 26 375
rect 17 371 26 373
rect 28 371 33 392
rect 35 384 40 392
rect 55 389 62 394
rect 55 387 57 389
rect 59 387 62 389
rect 55 385 62 387
rect 35 382 42 384
rect 35 380 38 382
rect 40 380 42 382
rect 57 380 62 385
rect 64 391 70 398
rect 103 396 110 398
rect 103 394 105 396
rect 107 394 110 396
rect 103 392 110 394
rect 64 384 72 391
rect 64 382 67 384
rect 69 382 72 384
rect 64 380 72 382
rect 35 378 42 380
rect 35 371 40 378
rect 66 378 72 380
rect 74 389 82 391
rect 74 387 77 389
rect 79 387 82 389
rect 74 382 82 387
rect 74 380 77 382
rect 79 380 82 382
rect 74 378 82 380
rect 84 382 91 391
rect 84 380 87 382
rect 89 380 91 382
rect 84 378 91 380
rect 105 371 110 392
rect 112 382 126 398
rect 112 380 115 382
rect 117 380 126 382
rect 128 396 136 398
rect 128 394 131 396
rect 133 394 136 396
rect 128 389 136 394
rect 128 387 131 389
rect 133 387 136 389
rect 128 380 136 387
rect 138 389 146 398
rect 138 387 141 389
rect 143 387 146 389
rect 138 380 146 387
rect 112 375 124 380
rect 112 373 115 375
rect 117 373 124 375
rect 112 371 124 373
rect 141 371 146 380
rect 148 383 153 398
rect 169 396 176 398
rect 169 394 171 396
rect 173 394 176 396
rect 169 389 176 394
rect 169 387 171 389
rect 173 387 176 389
rect 169 385 176 387
rect 148 381 155 383
rect 148 379 151 381
rect 153 379 155 381
rect 171 380 176 385
rect 178 391 184 398
rect 217 396 224 398
rect 217 394 219 396
rect 221 394 224 396
rect 217 392 224 394
rect 178 384 186 391
rect 178 382 181 384
rect 183 382 186 384
rect 178 380 186 382
rect 148 377 155 379
rect 148 371 153 377
rect 180 378 186 380
rect 188 389 196 391
rect 188 387 191 389
rect 193 387 196 389
rect 188 382 196 387
rect 188 380 191 382
rect 193 380 196 382
rect 188 378 196 380
rect 198 382 205 391
rect 198 380 201 382
rect 203 380 205 382
rect 198 378 205 380
rect 219 371 224 392
rect 226 382 240 398
rect 226 380 229 382
rect 231 380 240 382
rect 242 396 250 398
rect 242 394 245 396
rect 247 394 250 396
rect 242 389 250 394
rect 242 387 245 389
rect 247 387 250 389
rect 242 380 250 387
rect 252 389 260 398
rect 252 387 255 389
rect 257 387 260 389
rect 252 380 260 387
rect 226 375 238 380
rect 226 373 229 375
rect 231 373 238 375
rect 226 371 238 373
rect 255 371 260 380
rect 262 383 267 398
rect 301 391 307 398
rect 262 381 269 383
rect 262 379 265 381
rect 267 379 269 381
rect 262 377 269 379
rect 280 382 287 391
rect 280 380 282 382
rect 284 380 287 382
rect 280 378 287 380
rect 289 389 297 391
rect 289 387 292 389
rect 294 387 297 389
rect 289 382 297 387
rect 289 380 292 382
rect 294 380 297 382
rect 289 378 297 380
rect 299 384 307 391
rect 299 382 302 384
rect 304 382 307 384
rect 299 380 307 382
rect 309 396 316 398
rect 309 394 312 396
rect 314 394 316 396
rect 309 389 316 394
rect 322 397 329 399
rect 322 395 324 397
rect 326 395 329 397
rect 322 393 329 395
rect 324 391 329 393
rect 331 391 337 399
rect 309 387 312 389
rect 314 387 316 389
rect 309 385 316 387
rect 333 387 337 391
rect 368 387 373 389
rect 309 380 314 385
rect 333 383 339 387
rect 299 378 305 380
rect 262 371 267 377
rect 332 375 339 383
rect 332 373 334 375
rect 336 373 339 375
rect 332 371 339 373
rect 341 371 346 387
rect 348 385 356 387
rect 348 383 351 385
rect 353 383 356 385
rect 348 371 356 383
rect 358 371 363 387
rect 365 375 373 387
rect 365 373 368 375
rect 370 373 373 375
rect 365 371 373 373
rect 375 384 380 389
rect 391 384 396 389
rect 375 382 382 384
rect 375 380 378 382
rect 380 380 382 382
rect 375 378 382 380
rect 389 382 396 384
rect 389 380 391 382
rect 393 380 396 382
rect 389 378 396 380
rect 375 371 380 378
rect 391 371 396 378
rect 398 387 403 389
rect 434 391 440 399
rect 442 397 449 399
rect 442 395 445 397
rect 447 395 449 397
rect 442 393 449 395
rect 442 391 447 393
rect 434 387 438 391
rect 398 375 406 387
rect 398 373 401 375
rect 403 373 406 375
rect 398 371 406 373
rect 408 371 413 387
rect 415 385 423 387
rect 415 383 418 385
rect 420 383 423 385
rect 415 371 423 383
rect 425 371 430 387
rect 432 383 438 387
rect 458 384 463 389
rect 432 375 439 383
rect 456 382 463 384
rect 456 380 458 382
rect 460 380 463 382
rect 456 378 463 380
rect 432 373 435 375
rect 437 373 439 375
rect 432 371 439 373
rect 458 371 463 378
rect 465 387 470 389
rect 501 391 507 399
rect 509 397 516 399
rect 509 395 512 397
rect 514 395 516 397
rect 509 393 516 395
rect 524 394 529 399
rect 509 391 514 393
rect 522 392 529 394
rect 501 387 505 391
rect 465 375 473 387
rect 465 373 468 375
rect 470 373 473 375
rect 465 371 473 373
rect 475 371 480 387
rect 482 385 490 387
rect 482 383 485 385
rect 487 383 490 385
rect 482 371 490 383
rect 492 371 497 387
rect 499 383 505 387
rect 522 390 524 392
rect 526 390 529 392
rect 499 375 506 383
rect 522 385 529 390
rect 522 383 524 385
rect 526 383 529 385
rect 522 381 529 383
rect 531 392 539 399
rect 531 381 542 392
rect 499 373 502 375
rect 504 373 506 375
rect 533 375 542 381
rect 499 371 506 373
rect 533 373 535 375
rect 537 373 542 375
rect 533 371 542 373
rect 544 371 549 392
rect 551 384 556 392
rect 551 382 558 384
rect 566 383 571 398
rect 551 380 554 382
rect 556 380 558 382
rect 551 378 558 380
rect 564 381 571 383
rect 564 379 566 381
rect 568 379 571 381
rect 551 371 556 378
rect 564 377 571 379
rect 566 371 571 377
rect 573 389 581 398
rect 573 387 576 389
rect 578 387 581 389
rect 573 380 581 387
rect 583 396 591 398
rect 583 394 586 396
rect 588 394 591 396
rect 583 389 591 394
rect 583 387 586 389
rect 588 387 591 389
rect 583 380 591 387
rect 593 382 607 398
rect 593 380 602 382
rect 604 380 607 382
rect 573 371 578 380
rect 595 375 607 380
rect 595 373 602 375
rect 604 373 607 375
rect 595 371 607 373
rect 609 396 616 398
rect 609 394 612 396
rect 614 394 616 396
rect 609 392 616 394
rect 609 371 614 392
rect 17 357 26 359
rect 17 355 19 357
rect 21 355 26 357
rect 17 349 26 355
rect 6 347 13 349
rect 6 345 8 347
rect 10 345 13 347
rect 6 340 13 345
rect 6 338 8 340
rect 10 338 13 340
rect 6 336 13 338
rect 8 331 13 336
rect 15 338 26 349
rect 28 338 33 359
rect 35 352 40 359
rect 35 350 42 352
rect 66 350 72 352
rect 35 348 38 350
rect 40 348 42 350
rect 35 346 42 348
rect 35 338 40 346
rect 57 345 62 350
rect 55 343 62 345
rect 55 341 57 343
rect 59 341 62 343
rect 15 331 23 338
rect 55 336 62 341
rect 55 334 57 336
rect 59 334 62 336
rect 55 332 62 334
rect 64 348 72 350
rect 64 346 67 348
rect 69 346 72 348
rect 64 339 72 346
rect 74 350 82 352
rect 74 348 77 350
rect 79 348 82 350
rect 74 343 82 348
rect 74 341 77 343
rect 79 341 82 343
rect 74 339 82 341
rect 84 350 91 352
rect 84 348 87 350
rect 89 348 91 350
rect 84 339 91 348
rect 64 332 70 339
rect 105 338 110 359
rect 103 336 110 338
rect 103 334 105 336
rect 107 334 110 336
rect 103 332 110 334
rect 112 357 124 359
rect 112 355 115 357
rect 117 355 124 357
rect 112 350 124 355
rect 141 350 146 359
rect 112 348 115 350
rect 117 348 126 350
rect 112 332 126 348
rect 128 343 136 350
rect 128 341 131 343
rect 133 341 136 343
rect 128 336 136 341
rect 128 334 131 336
rect 133 334 136 336
rect 128 332 136 334
rect 138 343 146 350
rect 138 341 141 343
rect 143 341 146 343
rect 138 332 146 341
rect 148 353 153 359
rect 148 351 155 353
rect 148 349 151 351
rect 153 349 155 351
rect 180 350 186 352
rect 148 347 155 349
rect 148 332 153 347
rect 171 345 176 350
rect 169 343 176 345
rect 169 341 171 343
rect 173 341 176 343
rect 169 336 176 341
rect 169 334 171 336
rect 173 334 176 336
rect 169 332 176 334
rect 178 348 186 350
rect 178 346 181 348
rect 183 346 186 348
rect 178 339 186 346
rect 188 350 196 352
rect 188 348 191 350
rect 193 348 196 350
rect 188 343 196 348
rect 188 341 191 343
rect 193 341 196 343
rect 188 339 196 341
rect 198 350 205 352
rect 198 348 201 350
rect 203 348 205 350
rect 198 339 205 348
rect 178 332 184 339
rect 219 338 224 359
rect 217 336 224 338
rect 217 334 219 336
rect 221 334 224 336
rect 217 332 224 334
rect 226 357 238 359
rect 226 355 229 357
rect 231 355 238 357
rect 226 350 238 355
rect 255 350 260 359
rect 226 348 229 350
rect 231 348 240 350
rect 226 332 240 348
rect 242 343 250 350
rect 242 341 245 343
rect 247 341 250 343
rect 242 336 250 341
rect 242 334 245 336
rect 247 334 250 336
rect 242 332 250 334
rect 252 343 260 350
rect 252 341 255 343
rect 257 341 260 343
rect 252 332 260 341
rect 262 353 267 359
rect 262 351 269 353
rect 332 357 339 359
rect 332 355 334 357
rect 336 355 339 357
rect 262 349 265 351
rect 267 349 269 351
rect 262 347 269 349
rect 280 350 287 352
rect 280 348 282 350
rect 284 348 287 350
rect 262 332 267 347
rect 280 339 287 348
rect 289 350 297 352
rect 289 348 292 350
rect 294 348 297 350
rect 289 343 297 348
rect 289 341 292 343
rect 294 341 297 343
rect 289 339 297 341
rect 299 350 305 352
rect 299 348 307 350
rect 299 346 302 348
rect 304 346 307 348
rect 299 339 307 346
rect 301 332 307 339
rect 309 345 314 350
rect 332 347 339 355
rect 309 343 316 345
rect 309 341 312 343
rect 314 341 316 343
rect 309 336 316 341
rect 333 343 339 347
rect 341 343 346 359
rect 348 347 356 359
rect 348 345 351 347
rect 353 345 356 347
rect 348 343 356 345
rect 358 343 363 359
rect 365 357 373 359
rect 365 355 368 357
rect 370 355 373 357
rect 365 343 373 355
rect 333 339 337 343
rect 324 337 329 339
rect 309 334 312 336
rect 314 334 316 336
rect 309 332 316 334
rect 322 335 329 337
rect 322 333 324 335
rect 326 333 329 335
rect 322 331 329 333
rect 331 331 337 339
rect 368 341 373 343
rect 375 352 380 359
rect 391 352 396 359
rect 375 350 382 352
rect 375 348 378 350
rect 380 348 382 350
rect 375 346 382 348
rect 389 350 396 352
rect 389 348 391 350
rect 393 348 396 350
rect 389 346 396 348
rect 375 341 380 346
rect 391 341 396 346
rect 398 357 406 359
rect 398 355 401 357
rect 403 355 406 357
rect 398 343 406 355
rect 408 343 413 359
rect 415 347 423 359
rect 415 345 418 347
rect 420 345 423 347
rect 415 343 423 345
rect 425 343 430 359
rect 432 357 439 359
rect 432 355 435 357
rect 437 355 439 357
rect 432 347 439 355
rect 458 352 463 359
rect 456 350 463 352
rect 456 348 458 350
rect 460 348 463 350
rect 432 343 438 347
rect 456 346 463 348
rect 398 341 403 343
rect 434 339 438 343
rect 458 341 463 346
rect 465 357 473 359
rect 465 355 468 357
rect 470 355 473 357
rect 465 343 473 355
rect 475 343 480 359
rect 482 347 490 359
rect 482 345 485 347
rect 487 345 490 347
rect 482 343 490 345
rect 492 343 497 359
rect 499 357 506 359
rect 499 355 502 357
rect 504 355 506 357
rect 533 357 542 359
rect 499 347 506 355
rect 533 355 535 357
rect 537 355 542 357
rect 533 349 542 355
rect 499 343 505 347
rect 465 341 470 343
rect 434 331 440 339
rect 442 337 447 339
rect 442 335 449 337
rect 442 333 445 335
rect 447 333 449 335
rect 442 331 449 333
rect 501 339 505 343
rect 522 347 529 349
rect 522 345 524 347
rect 526 345 529 347
rect 522 340 529 345
rect 501 331 507 339
rect 509 337 514 339
rect 522 338 524 340
rect 526 338 529 340
rect 509 335 516 337
rect 522 336 529 338
rect 509 333 512 335
rect 514 333 516 335
rect 509 331 516 333
rect 524 331 529 336
rect 531 338 542 349
rect 544 338 549 359
rect 551 352 556 359
rect 566 353 571 359
rect 551 350 558 352
rect 551 348 554 350
rect 556 348 558 350
rect 551 346 558 348
rect 564 351 571 353
rect 564 349 566 351
rect 568 349 571 351
rect 564 347 571 349
rect 551 338 556 346
rect 531 331 539 338
rect 566 332 571 347
rect 573 350 578 359
rect 595 357 607 359
rect 595 355 602 357
rect 604 355 607 357
rect 595 350 607 355
rect 573 343 581 350
rect 573 341 576 343
rect 578 341 581 343
rect 573 332 581 341
rect 583 343 591 350
rect 583 341 586 343
rect 588 341 591 343
rect 583 336 591 341
rect 583 334 586 336
rect 588 334 591 336
rect 583 332 591 334
rect 593 348 602 350
rect 604 348 607 350
rect 593 332 607 348
rect 609 338 614 359
rect 609 336 616 338
rect 609 334 612 336
rect 614 334 616 336
rect 609 332 616 334
rect 8 250 13 255
rect 6 248 13 250
rect 6 246 8 248
rect 10 246 13 248
rect 6 241 13 246
rect 6 239 8 241
rect 10 239 13 241
rect 6 237 13 239
rect 15 248 23 255
rect 55 252 62 254
rect 55 250 57 252
rect 59 250 62 252
rect 15 237 26 248
rect 17 231 26 237
rect 17 229 19 231
rect 21 229 26 231
rect 17 227 26 229
rect 28 227 33 248
rect 35 240 40 248
rect 55 245 62 250
rect 55 243 57 245
rect 59 243 62 245
rect 55 241 62 243
rect 35 238 42 240
rect 35 236 38 238
rect 40 236 42 238
rect 57 236 62 241
rect 64 247 70 254
rect 103 252 110 254
rect 103 250 105 252
rect 107 250 110 252
rect 103 248 110 250
rect 64 240 72 247
rect 64 238 67 240
rect 69 238 72 240
rect 64 236 72 238
rect 35 234 42 236
rect 35 227 40 234
rect 66 234 72 236
rect 74 245 82 247
rect 74 243 77 245
rect 79 243 82 245
rect 74 238 82 243
rect 74 236 77 238
rect 79 236 82 238
rect 74 234 82 236
rect 84 238 91 247
rect 84 236 87 238
rect 89 236 91 238
rect 84 234 91 236
rect 105 227 110 248
rect 112 238 126 254
rect 112 236 115 238
rect 117 236 126 238
rect 128 252 136 254
rect 128 250 131 252
rect 133 250 136 252
rect 128 245 136 250
rect 128 243 131 245
rect 133 243 136 245
rect 128 236 136 243
rect 138 245 146 254
rect 138 243 141 245
rect 143 243 146 245
rect 138 236 146 243
rect 112 231 124 236
rect 112 229 115 231
rect 117 229 124 231
rect 112 227 124 229
rect 141 227 146 236
rect 148 239 153 254
rect 169 252 176 254
rect 169 250 171 252
rect 173 250 176 252
rect 169 245 176 250
rect 169 243 171 245
rect 173 243 176 245
rect 169 241 176 243
rect 148 237 155 239
rect 148 235 151 237
rect 153 235 155 237
rect 171 236 176 241
rect 178 247 184 254
rect 217 252 224 254
rect 217 250 219 252
rect 221 250 224 252
rect 217 248 224 250
rect 178 240 186 247
rect 178 238 181 240
rect 183 238 186 240
rect 178 236 186 238
rect 148 233 155 235
rect 148 227 153 233
rect 180 234 186 236
rect 188 245 196 247
rect 188 243 191 245
rect 193 243 196 245
rect 188 238 196 243
rect 188 236 191 238
rect 193 236 196 238
rect 188 234 196 236
rect 198 238 205 247
rect 198 236 201 238
rect 203 236 205 238
rect 198 234 205 236
rect 219 227 224 248
rect 226 238 240 254
rect 226 236 229 238
rect 231 236 240 238
rect 242 252 250 254
rect 242 250 245 252
rect 247 250 250 252
rect 242 245 250 250
rect 242 243 245 245
rect 247 243 250 245
rect 242 236 250 243
rect 252 245 260 254
rect 252 243 255 245
rect 257 243 260 245
rect 252 236 260 243
rect 226 231 238 236
rect 226 229 229 231
rect 231 229 238 231
rect 226 227 238 229
rect 255 227 260 236
rect 262 239 267 254
rect 301 247 307 254
rect 262 237 269 239
rect 262 235 265 237
rect 267 235 269 237
rect 262 233 269 235
rect 280 238 287 247
rect 280 236 282 238
rect 284 236 287 238
rect 280 234 287 236
rect 289 245 297 247
rect 289 243 292 245
rect 294 243 297 245
rect 289 238 297 243
rect 289 236 292 238
rect 294 236 297 238
rect 289 234 297 236
rect 299 240 307 247
rect 299 238 302 240
rect 304 238 307 240
rect 299 236 307 238
rect 309 252 316 254
rect 309 250 312 252
rect 314 250 316 252
rect 309 245 316 250
rect 322 253 329 255
rect 322 251 324 253
rect 326 251 329 253
rect 322 249 329 251
rect 324 247 329 249
rect 331 247 337 255
rect 309 243 312 245
rect 314 243 316 245
rect 309 241 316 243
rect 333 243 337 247
rect 368 243 373 245
rect 309 236 314 241
rect 333 239 339 243
rect 299 234 305 236
rect 262 227 267 233
rect 332 231 339 239
rect 332 229 334 231
rect 336 229 339 231
rect 332 227 339 229
rect 341 227 346 243
rect 348 241 356 243
rect 348 239 351 241
rect 353 239 356 241
rect 348 227 356 239
rect 358 227 363 243
rect 365 231 373 243
rect 365 229 368 231
rect 370 229 373 231
rect 365 227 373 229
rect 375 240 380 245
rect 391 240 396 245
rect 375 238 382 240
rect 375 236 378 238
rect 380 236 382 238
rect 375 234 382 236
rect 389 238 396 240
rect 389 236 391 238
rect 393 236 396 238
rect 389 234 396 236
rect 375 227 380 234
rect 391 227 396 234
rect 398 243 403 245
rect 434 247 440 255
rect 442 253 449 255
rect 442 251 445 253
rect 447 251 449 253
rect 442 249 449 251
rect 442 247 447 249
rect 434 243 438 247
rect 398 231 406 243
rect 398 229 401 231
rect 403 229 406 231
rect 398 227 406 229
rect 408 227 413 243
rect 415 241 423 243
rect 415 239 418 241
rect 420 239 423 241
rect 415 227 423 239
rect 425 227 430 243
rect 432 239 438 243
rect 458 240 463 245
rect 432 231 439 239
rect 456 238 463 240
rect 456 236 458 238
rect 460 236 463 238
rect 456 234 463 236
rect 432 229 435 231
rect 437 229 439 231
rect 432 227 439 229
rect 458 227 463 234
rect 465 243 470 245
rect 501 247 507 255
rect 509 253 516 255
rect 509 251 512 253
rect 514 251 516 253
rect 509 249 516 251
rect 524 250 529 255
rect 509 247 514 249
rect 522 248 529 250
rect 501 243 505 247
rect 465 231 473 243
rect 465 229 468 231
rect 470 229 473 231
rect 465 227 473 229
rect 475 227 480 243
rect 482 241 490 243
rect 482 239 485 241
rect 487 239 490 241
rect 482 227 490 239
rect 492 227 497 243
rect 499 239 505 243
rect 522 246 524 248
rect 526 246 529 248
rect 499 231 506 239
rect 522 241 529 246
rect 522 239 524 241
rect 526 239 529 241
rect 522 237 529 239
rect 531 248 539 255
rect 531 237 542 248
rect 499 229 502 231
rect 504 229 506 231
rect 533 231 542 237
rect 499 227 506 229
rect 533 229 535 231
rect 537 229 542 231
rect 533 227 542 229
rect 544 227 549 248
rect 551 240 556 248
rect 551 238 558 240
rect 566 239 571 254
rect 551 236 554 238
rect 556 236 558 238
rect 551 234 558 236
rect 564 237 571 239
rect 564 235 566 237
rect 568 235 571 237
rect 551 227 556 234
rect 564 233 571 235
rect 566 227 571 233
rect 573 245 581 254
rect 573 243 576 245
rect 578 243 581 245
rect 573 236 581 243
rect 583 252 591 254
rect 583 250 586 252
rect 588 250 591 252
rect 583 245 591 250
rect 583 243 586 245
rect 588 243 591 245
rect 583 236 591 243
rect 593 238 607 254
rect 593 236 602 238
rect 604 236 607 238
rect 573 227 578 236
rect 595 231 607 236
rect 595 229 602 231
rect 604 229 607 231
rect 595 227 607 229
rect 609 252 616 254
rect 609 250 612 252
rect 614 250 616 252
rect 609 248 616 250
rect 609 227 614 248
rect 17 213 26 215
rect 17 211 19 213
rect 21 211 26 213
rect 17 205 26 211
rect 6 203 13 205
rect 6 201 8 203
rect 10 201 13 203
rect 6 196 13 201
rect 6 194 8 196
rect 10 194 13 196
rect 6 192 13 194
rect 8 187 13 192
rect 15 194 26 205
rect 28 194 33 215
rect 35 208 40 215
rect 35 206 42 208
rect 66 206 72 208
rect 35 204 38 206
rect 40 204 42 206
rect 35 202 42 204
rect 35 194 40 202
rect 57 201 62 206
rect 55 199 62 201
rect 55 197 57 199
rect 59 197 62 199
rect 15 187 23 194
rect 55 192 62 197
rect 55 190 57 192
rect 59 190 62 192
rect 55 188 62 190
rect 64 204 72 206
rect 64 202 67 204
rect 69 202 72 204
rect 64 195 72 202
rect 74 206 82 208
rect 74 204 77 206
rect 79 204 82 206
rect 74 199 82 204
rect 74 197 77 199
rect 79 197 82 199
rect 74 195 82 197
rect 84 206 91 208
rect 84 204 87 206
rect 89 204 91 206
rect 84 195 91 204
rect 64 188 70 195
rect 105 194 110 215
rect 103 192 110 194
rect 103 190 105 192
rect 107 190 110 192
rect 103 188 110 190
rect 112 213 124 215
rect 112 211 115 213
rect 117 211 124 213
rect 112 206 124 211
rect 141 206 146 215
rect 112 204 115 206
rect 117 204 126 206
rect 112 188 126 204
rect 128 199 136 206
rect 128 197 131 199
rect 133 197 136 199
rect 128 192 136 197
rect 128 190 131 192
rect 133 190 136 192
rect 128 188 136 190
rect 138 199 146 206
rect 138 197 141 199
rect 143 197 146 199
rect 138 188 146 197
rect 148 209 153 215
rect 148 207 155 209
rect 148 205 151 207
rect 153 205 155 207
rect 180 206 186 208
rect 148 203 155 205
rect 148 188 153 203
rect 171 201 176 206
rect 169 199 176 201
rect 169 197 171 199
rect 173 197 176 199
rect 169 192 176 197
rect 169 190 171 192
rect 173 190 176 192
rect 169 188 176 190
rect 178 204 186 206
rect 178 202 181 204
rect 183 202 186 204
rect 178 195 186 202
rect 188 206 196 208
rect 188 204 191 206
rect 193 204 196 206
rect 188 199 196 204
rect 188 197 191 199
rect 193 197 196 199
rect 188 195 196 197
rect 198 206 205 208
rect 198 204 201 206
rect 203 204 205 206
rect 198 195 205 204
rect 178 188 184 195
rect 219 194 224 215
rect 217 192 224 194
rect 217 190 219 192
rect 221 190 224 192
rect 217 188 224 190
rect 226 213 238 215
rect 226 211 229 213
rect 231 211 238 213
rect 226 206 238 211
rect 255 206 260 215
rect 226 204 229 206
rect 231 204 240 206
rect 226 188 240 204
rect 242 199 250 206
rect 242 197 245 199
rect 247 197 250 199
rect 242 192 250 197
rect 242 190 245 192
rect 247 190 250 192
rect 242 188 250 190
rect 252 199 260 206
rect 252 197 255 199
rect 257 197 260 199
rect 252 188 260 197
rect 262 209 267 215
rect 262 207 269 209
rect 332 213 339 215
rect 332 211 334 213
rect 336 211 339 213
rect 262 205 265 207
rect 267 205 269 207
rect 262 203 269 205
rect 280 206 287 208
rect 280 204 282 206
rect 284 204 287 206
rect 262 188 267 203
rect 280 195 287 204
rect 289 206 297 208
rect 289 204 292 206
rect 294 204 297 206
rect 289 199 297 204
rect 289 197 292 199
rect 294 197 297 199
rect 289 195 297 197
rect 299 206 305 208
rect 299 204 307 206
rect 299 202 302 204
rect 304 202 307 204
rect 299 195 307 202
rect 301 188 307 195
rect 309 201 314 206
rect 332 203 339 211
rect 309 199 316 201
rect 309 197 312 199
rect 314 197 316 199
rect 309 192 316 197
rect 333 199 339 203
rect 341 199 346 215
rect 348 203 356 215
rect 348 201 351 203
rect 353 201 356 203
rect 348 199 356 201
rect 358 199 363 215
rect 365 213 373 215
rect 365 211 368 213
rect 370 211 373 213
rect 365 199 373 211
rect 333 195 337 199
rect 324 193 329 195
rect 309 190 312 192
rect 314 190 316 192
rect 309 188 316 190
rect 322 191 329 193
rect 322 189 324 191
rect 326 189 329 191
rect 322 187 329 189
rect 331 187 337 195
rect 368 197 373 199
rect 375 208 380 215
rect 391 208 396 215
rect 375 206 382 208
rect 375 204 378 206
rect 380 204 382 206
rect 375 202 382 204
rect 389 206 396 208
rect 389 204 391 206
rect 393 204 396 206
rect 389 202 396 204
rect 375 197 380 202
rect 391 197 396 202
rect 398 213 406 215
rect 398 211 401 213
rect 403 211 406 213
rect 398 199 406 211
rect 408 199 413 215
rect 415 203 423 215
rect 415 201 418 203
rect 420 201 423 203
rect 415 199 423 201
rect 425 199 430 215
rect 432 213 439 215
rect 432 211 435 213
rect 437 211 439 213
rect 432 203 439 211
rect 458 208 463 215
rect 456 206 463 208
rect 456 204 458 206
rect 460 204 463 206
rect 432 199 438 203
rect 456 202 463 204
rect 398 197 403 199
rect 434 195 438 199
rect 458 197 463 202
rect 465 213 473 215
rect 465 211 468 213
rect 470 211 473 213
rect 465 199 473 211
rect 475 199 480 215
rect 482 203 490 215
rect 482 201 485 203
rect 487 201 490 203
rect 482 199 490 201
rect 492 199 497 215
rect 499 213 506 215
rect 499 211 502 213
rect 504 211 506 213
rect 533 213 542 215
rect 499 203 506 211
rect 533 211 535 213
rect 537 211 542 213
rect 533 205 542 211
rect 499 199 505 203
rect 465 197 470 199
rect 434 187 440 195
rect 442 193 447 195
rect 442 191 449 193
rect 442 189 445 191
rect 447 189 449 191
rect 442 187 449 189
rect 501 195 505 199
rect 522 203 529 205
rect 522 201 524 203
rect 526 201 529 203
rect 522 196 529 201
rect 501 187 507 195
rect 509 193 514 195
rect 522 194 524 196
rect 526 194 529 196
rect 509 191 516 193
rect 522 192 529 194
rect 509 189 512 191
rect 514 189 516 191
rect 509 187 516 189
rect 524 187 529 192
rect 531 194 542 205
rect 544 194 549 215
rect 551 208 556 215
rect 566 209 571 215
rect 551 206 558 208
rect 551 204 554 206
rect 556 204 558 206
rect 551 202 558 204
rect 564 207 571 209
rect 564 205 566 207
rect 568 205 571 207
rect 564 203 571 205
rect 551 194 556 202
rect 531 187 539 194
rect 566 188 571 203
rect 573 206 578 215
rect 595 213 607 215
rect 595 211 602 213
rect 604 211 607 213
rect 595 206 607 211
rect 573 199 581 206
rect 573 197 576 199
rect 578 197 581 199
rect 573 188 581 197
rect 583 199 591 206
rect 583 197 586 199
rect 588 197 591 199
rect 583 192 591 197
rect 583 190 586 192
rect 588 190 591 192
rect 583 188 591 190
rect 593 204 602 206
rect 604 204 607 206
rect 593 188 607 204
rect 609 194 614 215
rect 609 192 616 194
rect 609 190 612 192
rect 614 190 616 192
rect 609 188 616 190
rect 8 106 13 111
rect 6 104 13 106
rect 6 102 8 104
rect 10 102 13 104
rect 6 97 13 102
rect 6 95 8 97
rect 10 95 13 97
rect 6 93 13 95
rect 15 104 23 111
rect 55 108 62 110
rect 55 106 57 108
rect 59 106 62 108
rect 15 93 26 104
rect 17 87 26 93
rect 17 85 19 87
rect 21 85 26 87
rect 17 83 26 85
rect 28 83 33 104
rect 35 96 40 104
rect 55 101 62 106
rect 55 99 57 101
rect 59 99 62 101
rect 55 97 62 99
rect 35 94 42 96
rect 35 92 38 94
rect 40 92 42 94
rect 57 92 62 97
rect 64 103 70 110
rect 103 108 110 110
rect 103 106 105 108
rect 107 106 110 108
rect 103 104 110 106
rect 64 96 72 103
rect 64 94 67 96
rect 69 94 72 96
rect 64 92 72 94
rect 35 90 42 92
rect 35 83 40 90
rect 66 90 72 92
rect 74 101 82 103
rect 74 99 77 101
rect 79 99 82 101
rect 74 94 82 99
rect 74 92 77 94
rect 79 92 82 94
rect 74 90 82 92
rect 84 94 91 103
rect 84 92 87 94
rect 89 92 91 94
rect 84 90 91 92
rect 105 83 110 104
rect 112 94 126 110
rect 112 92 115 94
rect 117 92 126 94
rect 128 108 136 110
rect 128 106 131 108
rect 133 106 136 108
rect 128 101 136 106
rect 128 99 131 101
rect 133 99 136 101
rect 128 92 136 99
rect 138 101 146 110
rect 138 99 141 101
rect 143 99 146 101
rect 138 92 146 99
rect 112 87 124 92
rect 112 85 115 87
rect 117 85 124 87
rect 112 83 124 85
rect 141 83 146 92
rect 148 95 153 110
rect 169 108 176 110
rect 169 106 171 108
rect 173 106 176 108
rect 169 101 176 106
rect 169 99 171 101
rect 173 99 176 101
rect 169 97 176 99
rect 148 93 155 95
rect 148 91 151 93
rect 153 91 155 93
rect 171 92 176 97
rect 178 103 184 110
rect 217 108 224 110
rect 217 106 219 108
rect 221 106 224 108
rect 217 104 224 106
rect 178 96 186 103
rect 178 94 181 96
rect 183 94 186 96
rect 178 92 186 94
rect 148 89 155 91
rect 148 83 153 89
rect 180 90 186 92
rect 188 101 196 103
rect 188 99 191 101
rect 193 99 196 101
rect 188 94 196 99
rect 188 92 191 94
rect 193 92 196 94
rect 188 90 196 92
rect 198 94 205 103
rect 198 92 201 94
rect 203 92 205 94
rect 198 90 205 92
rect 219 83 224 104
rect 226 94 240 110
rect 226 92 229 94
rect 231 92 240 94
rect 242 108 250 110
rect 242 106 245 108
rect 247 106 250 108
rect 242 101 250 106
rect 242 99 245 101
rect 247 99 250 101
rect 242 92 250 99
rect 252 101 260 110
rect 252 99 255 101
rect 257 99 260 101
rect 252 92 260 99
rect 226 87 238 92
rect 226 85 229 87
rect 231 85 238 87
rect 226 83 238 85
rect 255 83 260 92
rect 262 95 267 110
rect 301 103 307 110
rect 262 93 269 95
rect 262 91 265 93
rect 267 91 269 93
rect 262 89 269 91
rect 280 94 287 103
rect 280 92 282 94
rect 284 92 287 94
rect 280 90 287 92
rect 289 101 297 103
rect 289 99 292 101
rect 294 99 297 101
rect 289 94 297 99
rect 289 92 292 94
rect 294 92 297 94
rect 289 90 297 92
rect 299 96 307 103
rect 299 94 302 96
rect 304 94 307 96
rect 299 92 307 94
rect 309 108 316 110
rect 309 106 312 108
rect 314 106 316 108
rect 309 101 316 106
rect 322 109 329 111
rect 322 107 324 109
rect 326 107 329 109
rect 322 105 329 107
rect 324 103 329 105
rect 331 103 337 111
rect 309 99 312 101
rect 314 99 316 101
rect 309 97 316 99
rect 333 99 337 103
rect 368 99 373 101
rect 309 92 314 97
rect 333 95 339 99
rect 299 90 305 92
rect 262 83 267 89
rect 332 87 339 95
rect 332 85 334 87
rect 336 85 339 87
rect 332 83 339 85
rect 341 83 346 99
rect 348 97 356 99
rect 348 95 351 97
rect 353 95 356 97
rect 348 83 356 95
rect 358 83 363 99
rect 365 87 373 99
rect 365 85 368 87
rect 370 85 373 87
rect 365 83 373 85
rect 375 96 380 101
rect 391 96 396 101
rect 375 94 382 96
rect 375 92 378 94
rect 380 92 382 94
rect 375 90 382 92
rect 389 94 396 96
rect 389 92 391 94
rect 393 92 396 94
rect 389 90 396 92
rect 375 83 380 90
rect 391 83 396 90
rect 398 99 403 101
rect 434 103 440 111
rect 442 109 449 111
rect 442 107 445 109
rect 447 107 449 109
rect 442 105 449 107
rect 442 103 447 105
rect 434 99 438 103
rect 398 87 406 99
rect 398 85 401 87
rect 403 85 406 87
rect 398 83 406 85
rect 408 83 413 99
rect 415 97 423 99
rect 415 95 418 97
rect 420 95 423 97
rect 415 83 423 95
rect 425 83 430 99
rect 432 95 438 99
rect 458 96 463 101
rect 432 87 439 95
rect 456 94 463 96
rect 456 92 458 94
rect 460 92 463 94
rect 456 90 463 92
rect 432 85 435 87
rect 437 85 439 87
rect 432 83 439 85
rect 458 83 463 90
rect 465 99 470 101
rect 501 103 507 111
rect 509 109 516 111
rect 509 107 512 109
rect 514 107 516 109
rect 509 105 516 107
rect 524 106 529 111
rect 509 103 514 105
rect 522 104 529 106
rect 501 99 505 103
rect 465 87 473 99
rect 465 85 468 87
rect 470 85 473 87
rect 465 83 473 85
rect 475 83 480 99
rect 482 97 490 99
rect 482 95 485 97
rect 487 95 490 97
rect 482 83 490 95
rect 492 83 497 99
rect 499 95 505 99
rect 522 102 524 104
rect 526 102 529 104
rect 499 87 506 95
rect 522 97 529 102
rect 522 95 524 97
rect 526 95 529 97
rect 522 93 529 95
rect 531 104 539 111
rect 531 93 542 104
rect 499 85 502 87
rect 504 85 506 87
rect 533 87 542 93
rect 499 83 506 85
rect 533 85 535 87
rect 537 85 542 87
rect 533 83 542 85
rect 544 83 549 104
rect 551 96 556 104
rect 551 94 558 96
rect 566 95 571 110
rect 551 92 554 94
rect 556 92 558 94
rect 551 90 558 92
rect 564 93 571 95
rect 564 91 566 93
rect 568 91 571 93
rect 551 83 556 90
rect 564 89 571 91
rect 566 83 571 89
rect 573 101 581 110
rect 573 99 576 101
rect 578 99 581 101
rect 573 92 581 99
rect 583 108 591 110
rect 583 106 586 108
rect 588 106 591 108
rect 583 101 591 106
rect 583 99 586 101
rect 588 99 591 101
rect 583 92 591 99
rect 593 94 607 110
rect 593 92 602 94
rect 604 92 607 94
rect 573 83 578 92
rect 595 87 607 92
rect 595 85 602 87
rect 604 85 607 87
rect 595 83 607 85
rect 609 108 616 110
rect 609 106 612 108
rect 614 106 616 108
rect 609 104 616 106
rect 609 83 614 104
rect 17 69 26 71
rect 17 67 19 69
rect 21 67 26 69
rect 17 61 26 67
rect 6 59 13 61
rect 6 57 8 59
rect 10 57 13 59
rect 6 52 13 57
rect 6 50 8 52
rect 10 50 13 52
rect 6 48 13 50
rect 8 43 13 48
rect 15 50 26 61
rect 28 50 33 71
rect 35 64 40 71
rect 35 62 42 64
rect 66 62 72 64
rect 35 60 38 62
rect 40 60 42 62
rect 35 58 42 60
rect 35 50 40 58
rect 57 57 62 62
rect 55 55 62 57
rect 55 53 57 55
rect 59 53 62 55
rect 15 43 23 50
rect 55 48 62 53
rect 55 46 57 48
rect 59 46 62 48
rect 55 44 62 46
rect 64 60 72 62
rect 64 58 67 60
rect 69 58 72 60
rect 64 51 72 58
rect 74 62 82 64
rect 74 60 77 62
rect 79 60 82 62
rect 74 55 82 60
rect 74 53 77 55
rect 79 53 82 55
rect 74 51 82 53
rect 84 62 91 64
rect 84 60 87 62
rect 89 60 91 62
rect 84 51 91 60
rect 64 44 70 51
rect 105 50 110 71
rect 103 48 110 50
rect 103 46 105 48
rect 107 46 110 48
rect 103 44 110 46
rect 112 69 124 71
rect 112 67 115 69
rect 117 67 124 69
rect 112 62 124 67
rect 141 62 146 71
rect 112 60 115 62
rect 117 60 126 62
rect 112 44 126 60
rect 128 55 136 62
rect 128 53 131 55
rect 133 53 136 55
rect 128 48 136 53
rect 128 46 131 48
rect 133 46 136 48
rect 128 44 136 46
rect 138 55 146 62
rect 138 53 141 55
rect 143 53 146 55
rect 138 44 146 53
rect 148 65 153 71
rect 148 63 155 65
rect 148 61 151 63
rect 153 61 155 63
rect 180 62 186 64
rect 148 59 155 61
rect 148 44 153 59
rect 171 57 176 62
rect 169 55 176 57
rect 169 53 171 55
rect 173 53 176 55
rect 169 48 176 53
rect 169 46 171 48
rect 173 46 176 48
rect 169 44 176 46
rect 178 60 186 62
rect 178 58 181 60
rect 183 58 186 60
rect 178 51 186 58
rect 188 62 196 64
rect 188 60 191 62
rect 193 60 196 62
rect 188 55 196 60
rect 188 53 191 55
rect 193 53 196 55
rect 188 51 196 53
rect 198 62 205 64
rect 198 60 201 62
rect 203 60 205 62
rect 198 51 205 60
rect 178 44 184 51
rect 219 50 224 71
rect 217 48 224 50
rect 217 46 219 48
rect 221 46 224 48
rect 217 44 224 46
rect 226 69 238 71
rect 226 67 229 69
rect 231 67 238 69
rect 226 62 238 67
rect 255 62 260 71
rect 226 60 229 62
rect 231 60 240 62
rect 226 44 240 60
rect 242 55 250 62
rect 242 53 245 55
rect 247 53 250 55
rect 242 48 250 53
rect 242 46 245 48
rect 247 46 250 48
rect 242 44 250 46
rect 252 55 260 62
rect 252 53 255 55
rect 257 53 260 55
rect 252 44 260 53
rect 262 65 267 71
rect 262 63 269 65
rect 332 69 339 71
rect 332 67 334 69
rect 336 67 339 69
rect 262 61 265 63
rect 267 61 269 63
rect 262 59 269 61
rect 280 62 287 64
rect 280 60 282 62
rect 284 60 287 62
rect 262 44 267 59
rect 280 51 287 60
rect 289 62 297 64
rect 289 60 292 62
rect 294 60 297 62
rect 289 55 297 60
rect 289 53 292 55
rect 294 53 297 55
rect 289 51 297 53
rect 299 62 305 64
rect 299 60 307 62
rect 299 58 302 60
rect 304 58 307 60
rect 299 51 307 58
rect 301 44 307 51
rect 309 57 314 62
rect 332 59 339 67
rect 309 55 316 57
rect 309 53 312 55
rect 314 53 316 55
rect 309 48 316 53
rect 333 55 339 59
rect 341 55 346 71
rect 348 59 356 71
rect 348 57 351 59
rect 353 57 356 59
rect 348 55 356 57
rect 358 55 363 71
rect 365 69 373 71
rect 365 67 368 69
rect 370 67 373 69
rect 365 55 373 67
rect 333 51 337 55
rect 324 49 329 51
rect 309 46 312 48
rect 314 46 316 48
rect 309 44 316 46
rect 322 47 329 49
rect 322 45 324 47
rect 326 45 329 47
rect 322 43 329 45
rect 331 43 337 51
rect 368 53 373 55
rect 375 64 380 71
rect 391 64 396 71
rect 375 62 382 64
rect 375 60 378 62
rect 380 60 382 62
rect 375 58 382 60
rect 389 62 396 64
rect 389 60 391 62
rect 393 60 396 62
rect 389 58 396 60
rect 375 53 380 58
rect 391 53 396 58
rect 398 69 406 71
rect 398 67 401 69
rect 403 67 406 69
rect 398 55 406 67
rect 408 55 413 71
rect 415 59 423 71
rect 415 57 418 59
rect 420 57 423 59
rect 415 55 423 57
rect 425 55 430 71
rect 432 69 439 71
rect 432 67 435 69
rect 437 67 439 69
rect 432 59 439 67
rect 458 64 463 71
rect 456 62 463 64
rect 456 60 458 62
rect 460 60 463 62
rect 432 55 438 59
rect 456 58 463 60
rect 398 53 403 55
rect 434 51 438 55
rect 458 53 463 58
rect 465 69 473 71
rect 465 67 468 69
rect 470 67 473 69
rect 465 55 473 67
rect 475 55 480 71
rect 482 59 490 71
rect 482 57 485 59
rect 487 57 490 59
rect 482 55 490 57
rect 492 55 497 71
rect 499 69 506 71
rect 499 67 502 69
rect 504 67 506 69
rect 533 69 542 71
rect 499 59 506 67
rect 533 67 535 69
rect 537 67 542 69
rect 533 61 542 67
rect 499 55 505 59
rect 465 53 470 55
rect 434 43 440 51
rect 442 49 447 51
rect 442 47 449 49
rect 442 45 445 47
rect 447 45 449 47
rect 442 43 449 45
rect 501 51 505 55
rect 522 59 529 61
rect 522 57 524 59
rect 526 57 529 59
rect 522 52 529 57
rect 501 43 507 51
rect 509 49 514 51
rect 522 50 524 52
rect 526 50 529 52
rect 509 47 516 49
rect 522 48 529 50
rect 509 45 512 47
rect 514 45 516 47
rect 509 43 516 45
rect 524 43 529 48
rect 531 50 542 61
rect 544 50 549 71
rect 551 64 556 71
rect 566 65 571 71
rect 551 62 558 64
rect 551 60 554 62
rect 556 60 558 62
rect 551 58 558 60
rect 564 63 571 65
rect 564 61 566 63
rect 568 61 571 63
rect 564 59 571 61
rect 551 50 556 58
rect 531 43 539 50
rect 566 44 571 59
rect 573 62 578 71
rect 595 69 607 71
rect 595 67 602 69
rect 604 67 607 69
rect 595 62 607 67
rect 573 55 581 62
rect 573 53 576 55
rect 578 53 581 55
rect 573 44 581 53
rect 583 55 591 62
rect 583 53 586 55
rect 588 53 591 55
rect 583 48 591 53
rect 583 46 586 48
rect 588 46 591 48
rect 583 44 591 46
rect 593 60 602 62
rect 604 60 607 62
rect 593 44 607 60
rect 609 50 614 71
rect 609 48 616 50
rect 609 46 612 48
rect 614 46 616 48
rect 609 44 616 46
<< alu1 >>
rect 2 576 632 581
rect 2 574 9 576
rect 11 574 58 576
rect 60 574 68 576
rect 70 574 98 576
rect 100 574 151 576
rect 153 574 172 576
rect 174 574 182 576
rect 184 574 212 576
rect 214 574 265 576
rect 267 574 301 576
rect 303 574 311 576
rect 313 574 525 576
rect 527 574 566 576
rect 568 574 619 576
rect 621 574 632 576
rect 2 573 632 574
rect 55 564 67 568
rect 55 562 57 564
rect 59 562 67 564
rect 131 566 155 567
rect 6 559 11 561
rect 6 557 8 559
rect 10 557 11 559
rect 6 555 11 557
rect 6 536 10 555
rect 38 551 42 560
rect 6 534 8 536
rect 6 529 10 534
rect 6 527 8 529
rect 21 550 42 551
rect 21 548 25 550
rect 27 548 39 550
rect 41 548 42 550
rect 21 547 42 548
rect 21 541 35 543
rect 37 541 42 543
rect 21 539 42 541
rect 38 537 42 539
rect 55 542 59 562
rect 131 564 133 566
rect 135 564 155 566
rect 131 563 155 564
rect 79 559 84 560
rect 79 557 80 559
rect 82 557 84 559
rect 79 551 84 557
rect 55 540 60 542
rect 55 538 57 540
rect 59 538 60 540
rect 55 537 60 538
rect 38 533 60 537
rect 38 530 42 533
rect 55 531 57 533
rect 59 531 60 533
rect 70 550 84 551
rect 70 548 74 550
rect 76 548 84 550
rect 70 547 84 548
rect 103 559 116 560
rect 103 557 105 559
rect 107 557 116 559
rect 103 555 116 557
rect 103 554 113 555
rect 111 553 113 554
rect 115 553 116 555
rect 78 542 91 543
rect 78 540 84 542
rect 86 540 91 542
rect 78 539 91 540
rect 55 529 60 531
rect 6 523 19 527
rect 6 522 10 523
rect 87 535 91 539
rect 87 533 88 535
rect 90 533 91 535
rect 87 530 91 533
rect 95 542 100 544
rect 95 540 97 542
rect 99 540 100 542
rect 95 535 100 540
rect 111 546 116 553
rect 151 558 155 563
rect 151 556 152 558
rect 154 556 155 558
rect 95 533 97 535
rect 99 533 100 535
rect 95 528 100 533
rect 95 522 107 528
rect 151 535 155 556
rect 139 533 155 535
rect 139 531 141 533
rect 143 531 155 533
rect 139 530 155 531
rect 169 564 181 568
rect 169 562 171 564
rect 173 562 181 564
rect 245 566 269 567
rect 169 550 173 562
rect 245 564 247 566
rect 249 564 269 566
rect 245 563 269 564
rect 169 548 170 550
rect 172 548 173 550
rect 169 542 173 548
rect 193 559 198 560
rect 193 557 194 559
rect 196 557 198 559
rect 193 551 198 557
rect 169 540 174 542
rect 169 538 171 540
rect 173 538 174 540
rect 169 533 174 538
rect 169 531 171 533
rect 173 531 174 533
rect 184 550 198 551
rect 184 548 188 550
rect 190 548 198 550
rect 184 547 198 548
rect 217 559 230 560
rect 217 557 219 559
rect 221 557 230 559
rect 217 555 230 557
rect 217 554 227 555
rect 225 553 227 554
rect 229 553 230 555
rect 192 542 205 543
rect 192 540 198 542
rect 200 540 205 542
rect 192 539 205 540
rect 169 529 174 531
rect 201 535 205 539
rect 201 533 202 535
rect 204 533 205 535
rect 201 530 205 533
rect 209 542 214 544
rect 209 540 211 542
rect 213 540 214 542
rect 209 535 214 540
rect 225 546 230 553
rect 209 533 211 535
rect 213 533 214 535
rect 209 528 214 533
rect 209 522 221 528
rect 265 543 269 563
rect 287 551 292 560
rect 304 564 316 568
rect 304 562 312 564
rect 314 562 316 564
rect 287 550 301 551
rect 287 548 295 550
rect 297 548 301 550
rect 287 547 301 548
rect 265 541 266 543
rect 268 541 269 543
rect 265 535 269 541
rect 253 533 269 535
rect 253 531 255 533
rect 257 531 269 533
rect 253 530 269 531
rect 280 542 293 543
rect 280 540 285 542
rect 287 540 293 542
rect 280 539 293 540
rect 280 530 284 539
rect 312 558 316 562
rect 312 556 313 558
rect 315 556 316 558
rect 312 542 316 556
rect 311 540 316 542
rect 311 538 312 540
rect 314 538 316 540
rect 378 566 382 568
rect 377 564 382 566
rect 377 562 378 564
rect 380 562 382 564
rect 377 560 382 562
rect 329 558 342 559
rect 329 556 330 558
rect 332 556 342 558
rect 329 555 342 556
rect 336 550 342 555
rect 336 548 337 550
rect 339 548 342 550
rect 336 546 342 548
rect 362 545 366 552
rect 362 544 364 545
rect 354 543 364 544
rect 354 542 366 543
rect 354 540 355 542
rect 357 540 366 542
rect 354 538 366 540
rect 311 533 316 538
rect 311 531 312 533
rect 314 531 316 533
rect 311 529 316 531
rect 322 534 335 535
rect 322 532 332 534
rect 334 532 335 534
rect 322 531 335 532
rect 322 530 327 531
rect 378 550 382 560
rect 378 548 379 550
rect 381 548 382 550
rect 322 528 324 530
rect 326 528 327 530
rect 322 522 327 528
rect 378 527 382 548
rect 369 526 382 527
rect 369 524 378 526
rect 380 524 382 526
rect 369 523 382 524
rect 389 566 393 568
rect 389 564 394 566
rect 389 562 391 564
rect 393 562 394 564
rect 456 566 460 568
rect 389 560 394 562
rect 389 527 393 560
rect 429 558 442 559
rect 405 550 409 552
rect 405 548 406 550
rect 408 548 409 550
rect 405 545 409 548
rect 407 544 409 545
rect 407 543 417 544
rect 405 538 417 543
rect 429 556 437 558
rect 439 556 442 558
rect 429 555 442 556
rect 429 550 435 555
rect 429 548 432 550
rect 434 548 435 550
rect 429 546 435 548
rect 456 564 461 566
rect 456 562 458 564
rect 460 562 461 564
rect 564 566 588 567
rect 456 560 461 562
rect 456 558 460 560
rect 456 556 457 558
rect 459 556 460 558
rect 496 558 509 559
rect 436 531 449 535
rect 444 530 449 531
rect 389 526 402 527
rect 444 528 445 530
rect 447 528 449 530
rect 389 524 391 526
rect 393 524 402 526
rect 389 523 402 524
rect 444 522 449 528
rect 456 527 460 556
rect 472 545 476 552
rect 474 544 476 545
rect 474 543 484 544
rect 472 541 480 543
rect 482 541 484 543
rect 472 538 484 541
rect 496 556 505 558
rect 507 556 509 558
rect 496 555 509 556
rect 496 550 502 555
rect 496 548 499 550
rect 501 548 502 550
rect 496 546 502 548
rect 564 564 584 566
rect 586 564 588 566
rect 564 563 588 564
rect 522 559 527 561
rect 522 557 524 559
rect 526 557 527 559
rect 522 555 527 557
rect 522 542 526 555
rect 522 540 523 542
rect 525 540 526 542
rect 522 536 526 540
rect 554 551 558 560
rect 503 534 516 535
rect 503 532 504 534
rect 506 532 516 534
rect 503 531 516 532
rect 511 530 516 531
rect 456 526 469 527
rect 511 528 512 530
rect 514 528 516 530
rect 456 524 458 526
rect 460 524 469 526
rect 456 523 469 524
rect 511 522 516 528
rect 522 534 524 536
rect 522 529 526 534
rect 522 527 524 529
rect 537 550 558 551
rect 537 548 541 550
rect 543 548 558 550
rect 537 547 558 548
rect 564 558 568 563
rect 564 556 565 558
rect 567 556 568 558
rect 537 541 551 543
rect 553 541 558 543
rect 537 539 558 541
rect 554 530 558 539
rect 564 535 568 556
rect 603 555 616 560
rect 603 553 604 555
rect 606 554 616 555
rect 606 553 608 554
rect 564 533 580 535
rect 564 531 576 533
rect 578 531 580 533
rect 564 530 580 531
rect 603 546 608 553
rect 619 542 624 544
rect 619 540 620 542
rect 622 540 624 542
rect 522 523 535 527
rect 619 528 624 540
rect 522 522 526 523
rect 612 522 624 528
rect 2 516 632 517
rect 2 514 9 516
rect 11 514 58 516
rect 60 514 131 516
rect 133 514 172 516
rect 174 514 245 516
rect 247 514 311 516
rect 313 514 525 516
rect 527 514 586 516
rect 588 514 632 516
rect 2 504 632 514
rect 2 502 9 504
rect 11 502 58 504
rect 60 502 131 504
rect 133 502 172 504
rect 174 502 245 504
rect 247 502 311 504
rect 313 502 525 504
rect 527 502 586 504
rect 588 502 632 504
rect 2 501 632 502
rect 6 495 10 496
rect 6 491 19 495
rect 6 489 8 491
rect 6 484 10 489
rect 6 482 8 484
rect 6 463 10 482
rect 38 485 42 488
rect 55 487 60 489
rect 55 485 57 487
rect 59 485 60 487
rect 95 490 107 496
rect 38 481 60 485
rect 38 479 42 481
rect 21 477 42 479
rect 21 475 35 477
rect 37 475 42 477
rect 55 480 60 481
rect 55 478 57 480
rect 59 478 60 480
rect 55 476 60 478
rect 87 485 91 488
rect 87 483 88 485
rect 90 483 91 485
rect 6 461 11 463
rect 6 459 8 461
rect 10 459 11 461
rect 6 457 11 459
rect 21 470 42 471
rect 21 468 25 470
rect 27 468 39 470
rect 41 468 42 470
rect 21 467 42 468
rect 38 458 42 467
rect 55 456 59 476
rect 87 479 91 483
rect 78 478 91 479
rect 78 476 84 478
rect 86 476 91 478
rect 78 475 91 476
rect 95 485 100 490
rect 95 483 97 485
rect 99 483 100 485
rect 95 478 100 483
rect 95 476 97 478
rect 99 476 100 478
rect 95 474 100 476
rect 70 470 84 471
rect 70 468 74 470
rect 76 468 84 470
rect 70 467 84 468
rect 55 454 57 456
rect 59 454 67 456
rect 55 450 67 454
rect 79 461 84 467
rect 79 459 80 461
rect 82 459 84 461
rect 79 458 84 459
rect 111 465 116 472
rect 139 487 155 488
rect 139 485 141 487
rect 143 485 155 487
rect 139 483 155 485
rect 111 464 113 465
rect 103 463 113 464
rect 115 463 116 465
rect 103 461 116 463
rect 103 459 105 461
rect 107 459 116 461
rect 103 458 116 459
rect 151 462 155 483
rect 151 460 152 462
rect 154 460 155 462
rect 151 455 155 460
rect 131 454 155 455
rect 131 452 133 454
rect 135 452 155 454
rect 131 451 155 452
rect 169 487 174 489
rect 169 485 171 487
rect 173 485 174 487
rect 209 490 221 496
rect 169 480 174 485
rect 169 478 171 480
rect 173 478 174 480
rect 169 476 174 478
rect 201 485 205 488
rect 201 483 202 485
rect 204 483 205 485
rect 169 470 173 476
rect 169 468 170 470
rect 172 468 173 470
rect 169 456 173 468
rect 201 479 205 483
rect 192 478 205 479
rect 192 476 198 478
rect 200 476 205 478
rect 192 475 205 476
rect 209 485 214 490
rect 209 483 211 485
rect 213 483 214 485
rect 209 478 214 483
rect 209 476 211 478
rect 213 476 214 478
rect 209 474 214 476
rect 184 470 198 471
rect 184 468 188 470
rect 190 468 198 470
rect 184 467 198 468
rect 169 454 171 456
rect 173 454 181 456
rect 169 450 181 454
rect 193 461 198 467
rect 193 459 194 461
rect 196 459 198 461
rect 193 458 198 459
rect 225 465 230 472
rect 253 487 269 488
rect 253 485 255 487
rect 257 485 269 487
rect 253 483 269 485
rect 265 477 269 483
rect 265 475 266 477
rect 268 475 269 477
rect 280 479 284 488
rect 322 490 327 496
rect 369 494 382 495
rect 369 492 378 494
rect 380 492 382 494
rect 311 487 316 489
rect 280 478 293 479
rect 280 476 285 478
rect 287 476 293 478
rect 280 475 293 476
rect 225 464 227 465
rect 217 463 227 464
rect 229 463 230 465
rect 217 461 230 463
rect 217 459 219 461
rect 221 459 230 461
rect 217 458 230 459
rect 265 455 269 475
rect 287 470 301 471
rect 287 468 295 470
rect 297 468 301 470
rect 287 467 301 468
rect 311 485 312 487
rect 314 485 316 487
rect 311 480 316 485
rect 322 488 324 490
rect 326 488 327 490
rect 369 491 382 492
rect 322 487 327 488
rect 322 486 335 487
rect 322 484 332 486
rect 334 484 335 486
rect 322 483 335 484
rect 311 478 312 480
rect 314 478 316 480
rect 311 476 316 478
rect 287 458 292 467
rect 312 462 316 476
rect 312 460 313 462
rect 315 460 316 462
rect 312 456 316 460
rect 245 454 269 455
rect 245 452 247 454
rect 249 452 269 454
rect 245 451 269 452
rect 304 454 312 456
rect 314 454 316 456
rect 304 450 316 454
rect 336 470 342 472
rect 336 468 337 470
rect 339 468 342 470
rect 336 463 342 468
rect 329 462 342 463
rect 329 460 330 462
rect 332 460 342 462
rect 354 478 366 480
rect 354 476 355 478
rect 357 476 366 478
rect 354 475 366 476
rect 354 474 364 475
rect 362 473 364 474
rect 362 466 366 473
rect 378 470 382 491
rect 378 468 379 470
rect 381 468 382 470
rect 329 459 342 460
rect 378 458 382 468
rect 377 456 382 458
rect 377 454 378 456
rect 380 454 382 456
rect 377 452 382 454
rect 378 450 382 452
rect 389 494 402 495
rect 389 492 391 494
rect 393 492 402 494
rect 389 491 402 492
rect 389 458 393 491
rect 444 490 449 496
rect 444 488 445 490
rect 447 488 449 490
rect 444 487 449 488
rect 436 483 449 487
rect 456 494 469 495
rect 456 492 458 494
rect 460 492 469 494
rect 456 491 469 492
rect 405 475 417 480
rect 407 474 417 475
rect 407 473 409 474
rect 405 470 409 473
rect 405 468 406 470
rect 408 468 409 470
rect 405 466 409 468
rect 429 470 435 472
rect 429 468 432 470
rect 434 468 435 470
rect 429 463 435 468
rect 429 462 442 463
rect 429 460 437 462
rect 439 460 442 462
rect 429 459 442 460
rect 389 456 394 458
rect 389 454 391 456
rect 393 454 394 456
rect 389 452 394 454
rect 389 450 393 452
rect 456 462 460 491
rect 511 490 516 496
rect 511 488 512 490
rect 514 488 516 490
rect 511 487 516 488
rect 503 486 516 487
rect 503 484 504 486
rect 506 484 516 486
rect 503 483 516 484
rect 522 495 526 496
rect 522 491 535 495
rect 522 489 524 491
rect 522 484 526 489
rect 522 482 524 484
rect 472 477 484 480
rect 472 475 480 477
rect 482 475 484 477
rect 474 474 484 475
rect 474 473 476 474
rect 456 460 457 462
rect 459 460 460 462
rect 472 466 476 473
rect 456 458 460 460
rect 496 470 502 472
rect 496 468 499 470
rect 501 468 502 470
rect 496 463 502 468
rect 496 462 509 463
rect 496 460 505 462
rect 507 460 509 462
rect 496 459 509 460
rect 456 456 461 458
rect 456 454 458 456
rect 460 454 461 456
rect 456 452 461 454
rect 456 450 460 452
rect 522 478 526 482
rect 522 476 523 478
rect 525 476 526 478
rect 522 463 526 476
rect 554 479 558 488
rect 537 477 558 479
rect 537 475 551 477
rect 553 475 558 477
rect 564 487 580 488
rect 564 485 576 487
rect 578 485 580 487
rect 564 483 580 485
rect 522 461 527 463
rect 522 459 524 461
rect 526 459 527 461
rect 522 457 527 459
rect 537 470 558 471
rect 537 468 541 470
rect 543 468 558 470
rect 537 467 558 468
rect 554 458 558 467
rect 564 462 568 483
rect 612 490 624 496
rect 564 460 565 462
rect 567 460 568 462
rect 564 455 568 460
rect 603 465 608 472
rect 619 478 624 490
rect 619 476 620 478
rect 622 476 624 478
rect 619 474 624 476
rect 603 463 604 465
rect 606 464 608 465
rect 606 463 616 464
rect 603 458 616 463
rect 564 454 588 455
rect 564 452 584 454
rect 586 452 588 454
rect 564 451 588 452
rect 2 444 632 445
rect 2 442 9 444
rect 11 442 58 444
rect 60 442 68 444
rect 70 442 98 444
rect 100 442 151 444
rect 153 442 172 444
rect 174 442 182 444
rect 184 442 212 444
rect 214 442 265 444
rect 267 442 301 444
rect 303 442 311 444
rect 313 442 525 444
rect 527 442 566 444
rect 568 442 619 444
rect 621 442 632 444
rect 2 432 632 442
rect 2 430 9 432
rect 11 430 58 432
rect 60 430 68 432
rect 70 430 98 432
rect 100 430 151 432
rect 153 430 172 432
rect 174 430 182 432
rect 184 430 212 432
rect 214 430 265 432
rect 267 430 301 432
rect 303 430 311 432
rect 313 430 525 432
rect 527 430 566 432
rect 568 430 619 432
rect 621 430 632 432
rect 2 429 632 430
rect 55 420 67 424
rect 55 418 57 420
rect 59 418 67 420
rect 131 422 155 423
rect 6 415 11 417
rect 6 413 8 415
rect 10 413 11 415
rect 6 411 11 413
rect 6 392 10 411
rect 38 407 42 416
rect 6 390 8 392
rect 6 385 10 390
rect 6 383 8 385
rect 21 406 42 407
rect 21 404 25 406
rect 27 404 39 406
rect 41 404 42 406
rect 21 403 42 404
rect 21 397 35 399
rect 37 397 42 399
rect 21 395 42 397
rect 38 393 42 395
rect 55 398 59 418
rect 131 420 133 422
rect 135 420 155 422
rect 131 419 155 420
rect 79 415 84 416
rect 79 413 80 415
rect 82 413 84 415
rect 79 407 84 413
rect 55 396 60 398
rect 55 394 57 396
rect 59 394 60 396
rect 55 393 60 394
rect 38 389 60 393
rect 38 386 42 389
rect 55 387 57 389
rect 59 387 60 389
rect 70 406 84 407
rect 70 404 74 406
rect 76 404 84 406
rect 70 403 84 404
rect 103 415 116 416
rect 103 413 105 415
rect 107 413 116 415
rect 103 411 116 413
rect 103 410 113 411
rect 111 409 113 410
rect 115 409 116 411
rect 78 398 91 399
rect 78 396 84 398
rect 86 396 91 398
rect 78 395 91 396
rect 55 385 60 387
rect 6 379 19 383
rect 6 378 10 379
rect 87 391 91 395
rect 87 389 88 391
rect 90 389 91 391
rect 87 386 91 389
rect 95 398 100 400
rect 95 396 97 398
rect 99 396 100 398
rect 95 391 100 396
rect 111 402 116 409
rect 151 414 155 419
rect 151 412 152 414
rect 154 412 155 414
rect 95 389 97 391
rect 99 389 100 391
rect 95 384 100 389
rect 95 378 107 384
rect 151 391 155 412
rect 139 389 155 391
rect 139 387 141 389
rect 143 387 155 389
rect 139 386 155 387
rect 169 420 181 424
rect 169 418 171 420
rect 173 418 181 420
rect 245 422 269 423
rect 169 406 173 418
rect 245 420 247 422
rect 249 420 269 422
rect 245 419 269 420
rect 169 404 170 406
rect 172 404 173 406
rect 169 398 173 404
rect 193 415 198 416
rect 193 413 194 415
rect 196 413 198 415
rect 193 407 198 413
rect 169 396 174 398
rect 169 394 171 396
rect 173 394 174 396
rect 169 389 174 394
rect 169 387 171 389
rect 173 387 174 389
rect 184 406 198 407
rect 184 404 188 406
rect 190 404 198 406
rect 184 403 198 404
rect 217 415 230 416
rect 217 413 219 415
rect 221 413 230 415
rect 217 411 230 413
rect 217 410 227 411
rect 225 409 227 410
rect 229 409 230 411
rect 192 398 205 399
rect 192 396 198 398
rect 200 396 205 398
rect 192 395 205 396
rect 169 385 174 387
rect 201 391 205 395
rect 201 389 202 391
rect 204 389 205 391
rect 201 386 205 389
rect 209 398 214 400
rect 209 396 211 398
rect 213 396 214 398
rect 209 391 214 396
rect 225 402 230 409
rect 209 389 211 391
rect 213 389 214 391
rect 209 384 214 389
rect 209 378 221 384
rect 265 399 269 419
rect 287 407 292 416
rect 304 420 316 424
rect 304 418 312 420
rect 314 418 316 420
rect 287 406 301 407
rect 287 404 295 406
rect 297 404 301 406
rect 287 403 301 404
rect 265 397 266 399
rect 268 397 269 399
rect 265 391 269 397
rect 253 389 269 391
rect 253 387 255 389
rect 257 387 269 389
rect 253 386 269 387
rect 280 398 293 399
rect 280 396 285 398
rect 287 396 293 398
rect 280 395 293 396
rect 280 386 284 395
rect 312 414 316 418
rect 312 412 313 414
rect 315 412 316 414
rect 312 398 316 412
rect 311 396 316 398
rect 311 394 312 396
rect 314 394 316 396
rect 378 422 382 424
rect 377 420 382 422
rect 377 418 378 420
rect 380 418 382 420
rect 377 416 382 418
rect 329 414 342 415
rect 329 412 330 414
rect 332 412 342 414
rect 329 411 342 412
rect 336 406 342 411
rect 336 404 337 406
rect 339 404 342 406
rect 336 402 342 404
rect 362 401 366 408
rect 362 400 364 401
rect 354 399 364 400
rect 354 398 366 399
rect 354 396 355 398
rect 357 396 366 398
rect 354 394 366 396
rect 311 389 316 394
rect 311 387 312 389
rect 314 387 316 389
rect 311 385 316 387
rect 322 390 335 391
rect 322 388 332 390
rect 334 388 335 390
rect 322 387 335 388
rect 322 386 327 387
rect 378 406 382 416
rect 378 404 379 406
rect 381 404 382 406
rect 322 384 324 386
rect 326 384 327 386
rect 322 378 327 384
rect 378 383 382 404
rect 369 382 382 383
rect 369 380 378 382
rect 380 380 382 382
rect 369 379 382 380
rect 389 422 393 424
rect 389 420 394 422
rect 389 418 391 420
rect 393 418 394 420
rect 456 422 460 424
rect 389 416 394 418
rect 389 383 393 416
rect 429 414 442 415
rect 405 406 409 408
rect 405 404 406 406
rect 408 404 409 406
rect 405 401 409 404
rect 407 400 409 401
rect 407 399 417 400
rect 405 394 417 399
rect 429 412 437 414
rect 439 412 442 414
rect 429 411 442 412
rect 429 406 435 411
rect 429 404 432 406
rect 434 404 435 406
rect 429 402 435 404
rect 456 420 461 422
rect 456 418 458 420
rect 460 418 461 420
rect 564 422 588 423
rect 456 416 461 418
rect 456 414 460 416
rect 456 412 457 414
rect 459 412 460 414
rect 496 414 509 415
rect 436 387 449 391
rect 444 386 449 387
rect 389 382 402 383
rect 444 384 445 386
rect 447 384 449 386
rect 389 380 391 382
rect 393 380 402 382
rect 389 379 402 380
rect 444 378 449 384
rect 456 383 460 412
rect 472 401 476 408
rect 474 400 476 401
rect 474 399 484 400
rect 472 397 480 399
rect 482 397 484 399
rect 472 394 484 397
rect 496 412 505 414
rect 507 412 509 414
rect 496 411 509 412
rect 496 406 502 411
rect 496 404 499 406
rect 501 404 502 406
rect 496 402 502 404
rect 564 420 584 422
rect 586 420 588 422
rect 564 419 588 420
rect 522 415 527 417
rect 522 413 524 415
rect 526 413 527 415
rect 522 411 527 413
rect 522 398 526 411
rect 522 396 523 398
rect 525 396 526 398
rect 522 392 526 396
rect 554 407 558 416
rect 503 390 516 391
rect 503 388 504 390
rect 506 388 516 390
rect 503 387 516 388
rect 511 386 516 387
rect 456 382 469 383
rect 511 384 512 386
rect 514 384 516 386
rect 456 380 458 382
rect 460 380 469 382
rect 456 379 469 380
rect 511 378 516 384
rect 522 390 524 392
rect 522 385 526 390
rect 522 383 524 385
rect 537 406 558 407
rect 537 404 541 406
rect 543 404 558 406
rect 537 403 558 404
rect 564 414 568 419
rect 564 412 565 414
rect 567 412 568 414
rect 537 397 551 399
rect 553 397 558 399
rect 537 395 558 397
rect 554 386 558 395
rect 564 391 568 412
rect 603 411 616 416
rect 603 409 604 411
rect 606 410 616 411
rect 606 409 608 410
rect 564 389 580 391
rect 564 387 576 389
rect 578 387 580 389
rect 564 386 580 387
rect 603 402 608 409
rect 619 398 624 400
rect 619 396 620 398
rect 622 396 624 398
rect 522 379 535 383
rect 619 384 624 396
rect 522 378 526 379
rect 612 378 624 384
rect 2 372 632 373
rect 2 370 9 372
rect 11 370 58 372
rect 60 370 131 372
rect 133 370 172 372
rect 174 370 245 372
rect 247 370 311 372
rect 313 370 525 372
rect 527 370 586 372
rect 588 370 632 372
rect 2 360 632 370
rect 2 358 9 360
rect 11 358 58 360
rect 60 358 131 360
rect 133 358 172 360
rect 174 358 245 360
rect 247 358 311 360
rect 313 358 525 360
rect 527 358 586 360
rect 588 358 632 360
rect 2 357 632 358
rect 6 351 10 352
rect 6 347 19 351
rect 6 345 8 347
rect 6 340 10 345
rect 6 338 8 340
rect 6 319 10 338
rect 38 341 42 344
rect 55 343 60 345
rect 55 341 57 343
rect 59 341 60 343
rect 95 346 107 352
rect 38 337 60 341
rect 38 335 42 337
rect 21 333 42 335
rect 21 331 35 333
rect 37 331 42 333
rect 55 336 60 337
rect 55 334 57 336
rect 59 334 60 336
rect 55 332 60 334
rect 87 341 91 344
rect 87 339 88 341
rect 90 339 91 341
rect 6 317 11 319
rect 6 315 8 317
rect 10 315 11 317
rect 6 313 11 315
rect 21 326 42 327
rect 21 324 25 326
rect 27 324 39 326
rect 41 324 42 326
rect 21 323 42 324
rect 38 314 42 323
rect 55 312 59 332
rect 87 335 91 339
rect 78 334 91 335
rect 78 332 84 334
rect 86 332 91 334
rect 78 331 91 332
rect 95 341 100 346
rect 95 339 97 341
rect 99 339 100 341
rect 95 334 100 339
rect 95 332 97 334
rect 99 332 100 334
rect 95 330 100 332
rect 70 326 84 327
rect 70 324 74 326
rect 76 324 84 326
rect 70 323 84 324
rect 55 310 57 312
rect 59 310 67 312
rect 55 306 67 310
rect 79 317 84 323
rect 79 315 80 317
rect 82 315 84 317
rect 79 314 84 315
rect 111 321 116 328
rect 139 343 155 344
rect 139 341 141 343
rect 143 341 155 343
rect 139 339 155 341
rect 111 320 113 321
rect 103 319 113 320
rect 115 319 116 321
rect 103 317 116 319
rect 103 315 105 317
rect 107 315 116 317
rect 103 314 116 315
rect 151 318 155 339
rect 151 316 152 318
rect 154 316 155 318
rect 151 311 155 316
rect 131 310 155 311
rect 131 308 133 310
rect 135 308 155 310
rect 131 307 155 308
rect 169 343 174 345
rect 169 341 171 343
rect 173 341 174 343
rect 209 346 221 352
rect 169 336 174 341
rect 169 334 171 336
rect 173 334 174 336
rect 169 332 174 334
rect 201 341 205 344
rect 201 339 202 341
rect 204 339 205 341
rect 169 326 173 332
rect 169 324 170 326
rect 172 324 173 326
rect 169 312 173 324
rect 201 335 205 339
rect 192 334 205 335
rect 192 332 198 334
rect 200 332 205 334
rect 192 331 205 332
rect 209 341 214 346
rect 209 339 211 341
rect 213 339 214 341
rect 209 334 214 339
rect 209 332 211 334
rect 213 332 214 334
rect 209 330 214 332
rect 184 326 198 327
rect 184 324 188 326
rect 190 324 198 326
rect 184 323 198 324
rect 169 310 171 312
rect 173 310 181 312
rect 169 306 181 310
rect 193 317 198 323
rect 193 315 194 317
rect 196 315 198 317
rect 193 314 198 315
rect 225 321 230 328
rect 253 343 269 344
rect 253 341 255 343
rect 257 341 269 343
rect 253 339 269 341
rect 265 333 269 339
rect 265 331 266 333
rect 268 331 269 333
rect 280 335 284 344
rect 322 346 327 352
rect 369 350 382 351
rect 369 348 378 350
rect 380 348 382 350
rect 311 343 316 345
rect 280 334 293 335
rect 280 332 285 334
rect 287 332 293 334
rect 280 331 293 332
rect 225 320 227 321
rect 217 319 227 320
rect 229 319 230 321
rect 217 317 230 319
rect 217 315 219 317
rect 221 315 230 317
rect 217 314 230 315
rect 265 311 269 331
rect 287 326 301 327
rect 287 324 295 326
rect 297 324 301 326
rect 287 323 301 324
rect 311 341 312 343
rect 314 341 316 343
rect 311 336 316 341
rect 322 344 324 346
rect 326 344 327 346
rect 369 347 382 348
rect 322 343 327 344
rect 322 342 335 343
rect 322 340 332 342
rect 334 340 335 342
rect 322 339 335 340
rect 311 334 312 336
rect 314 334 316 336
rect 311 332 316 334
rect 287 314 292 323
rect 312 318 316 332
rect 312 316 313 318
rect 315 316 316 318
rect 312 312 316 316
rect 245 310 269 311
rect 245 308 247 310
rect 249 308 269 310
rect 245 307 269 308
rect 304 310 312 312
rect 314 310 316 312
rect 304 306 316 310
rect 336 326 342 328
rect 336 324 337 326
rect 339 324 342 326
rect 336 319 342 324
rect 329 318 342 319
rect 329 316 330 318
rect 332 316 342 318
rect 354 334 366 336
rect 354 332 355 334
rect 357 332 366 334
rect 354 331 366 332
rect 354 330 364 331
rect 362 329 364 330
rect 362 322 366 329
rect 378 326 382 347
rect 378 324 379 326
rect 381 324 382 326
rect 329 315 342 316
rect 378 314 382 324
rect 377 312 382 314
rect 377 310 378 312
rect 380 310 382 312
rect 377 308 382 310
rect 378 306 382 308
rect 389 350 402 351
rect 389 348 391 350
rect 393 348 402 350
rect 389 347 402 348
rect 389 314 393 347
rect 444 346 449 352
rect 444 344 445 346
rect 447 344 449 346
rect 444 343 449 344
rect 436 339 449 343
rect 456 350 469 351
rect 456 348 458 350
rect 460 348 469 350
rect 456 347 469 348
rect 405 331 417 336
rect 407 330 417 331
rect 407 329 409 330
rect 405 326 409 329
rect 405 324 406 326
rect 408 324 409 326
rect 405 322 409 324
rect 429 326 435 328
rect 429 324 432 326
rect 434 324 435 326
rect 429 319 435 324
rect 429 318 442 319
rect 429 316 437 318
rect 439 316 442 318
rect 429 315 442 316
rect 389 312 394 314
rect 389 310 391 312
rect 393 310 394 312
rect 389 308 394 310
rect 389 306 393 308
rect 456 318 460 347
rect 511 346 516 352
rect 511 344 512 346
rect 514 344 516 346
rect 511 343 516 344
rect 503 342 516 343
rect 503 340 504 342
rect 506 340 516 342
rect 503 339 516 340
rect 522 351 526 352
rect 522 347 535 351
rect 522 345 524 347
rect 522 340 526 345
rect 522 338 524 340
rect 472 333 484 336
rect 472 331 480 333
rect 482 331 484 333
rect 474 330 484 331
rect 474 329 476 330
rect 456 316 457 318
rect 459 316 460 318
rect 472 322 476 329
rect 456 314 460 316
rect 496 326 502 328
rect 496 324 499 326
rect 501 324 502 326
rect 496 319 502 324
rect 496 318 509 319
rect 496 316 505 318
rect 507 316 509 318
rect 496 315 509 316
rect 456 312 461 314
rect 456 310 458 312
rect 460 310 461 312
rect 456 308 461 310
rect 456 306 460 308
rect 522 334 526 338
rect 522 332 523 334
rect 525 332 526 334
rect 522 319 526 332
rect 554 335 558 344
rect 537 333 558 335
rect 537 331 551 333
rect 553 331 558 333
rect 564 343 580 344
rect 564 341 576 343
rect 578 341 580 343
rect 564 339 580 341
rect 522 317 527 319
rect 522 315 524 317
rect 526 315 527 317
rect 522 313 527 315
rect 537 326 558 327
rect 537 324 541 326
rect 543 324 558 326
rect 537 323 558 324
rect 554 314 558 323
rect 564 318 568 339
rect 612 346 624 352
rect 564 316 565 318
rect 567 316 568 318
rect 564 311 568 316
rect 603 321 608 328
rect 619 334 624 346
rect 619 332 620 334
rect 622 332 624 334
rect 619 330 624 332
rect 603 319 604 321
rect 606 320 608 321
rect 606 319 616 320
rect 603 314 616 319
rect 564 310 588 311
rect 564 308 584 310
rect 586 308 588 310
rect 564 307 588 308
rect 2 300 632 301
rect 2 298 9 300
rect 11 298 58 300
rect 60 298 68 300
rect 70 298 98 300
rect 100 298 151 300
rect 153 298 172 300
rect 174 298 182 300
rect 184 298 212 300
rect 214 298 265 300
rect 267 298 301 300
rect 303 298 311 300
rect 313 298 525 300
rect 527 298 566 300
rect 568 298 619 300
rect 621 298 632 300
rect 2 288 632 298
rect 2 286 9 288
rect 11 286 58 288
rect 60 286 68 288
rect 70 286 98 288
rect 100 286 151 288
rect 153 286 172 288
rect 174 286 182 288
rect 184 286 212 288
rect 214 286 265 288
rect 267 286 301 288
rect 303 286 311 288
rect 313 286 525 288
rect 527 286 566 288
rect 568 286 619 288
rect 621 286 632 288
rect 2 285 632 286
rect 55 276 67 280
rect 55 274 57 276
rect 59 274 67 276
rect 131 278 155 279
rect 6 271 11 273
rect 6 269 8 271
rect 10 269 11 271
rect 6 267 11 269
rect 6 248 10 267
rect 38 263 42 272
rect 6 246 8 248
rect 6 241 10 246
rect 6 239 8 241
rect 21 262 42 263
rect 21 260 25 262
rect 27 260 39 262
rect 41 260 42 262
rect 21 259 42 260
rect 21 253 35 255
rect 37 253 42 255
rect 21 251 42 253
rect 38 249 42 251
rect 55 254 59 274
rect 131 276 133 278
rect 135 276 155 278
rect 131 275 155 276
rect 79 271 84 272
rect 79 269 80 271
rect 82 269 84 271
rect 79 263 84 269
rect 55 252 60 254
rect 55 250 57 252
rect 59 250 60 252
rect 55 249 60 250
rect 38 245 60 249
rect 38 242 42 245
rect 55 243 57 245
rect 59 243 60 245
rect 70 262 84 263
rect 70 260 74 262
rect 76 260 84 262
rect 70 259 84 260
rect 103 271 116 272
rect 103 269 105 271
rect 107 269 116 271
rect 103 267 116 269
rect 103 266 113 267
rect 111 265 113 266
rect 115 265 116 267
rect 78 254 91 255
rect 78 252 84 254
rect 86 252 91 254
rect 78 251 91 252
rect 55 241 60 243
rect 6 235 19 239
rect 6 234 10 235
rect 87 247 91 251
rect 87 245 88 247
rect 90 245 91 247
rect 87 242 91 245
rect 95 254 100 256
rect 95 252 97 254
rect 99 252 100 254
rect 95 247 100 252
rect 111 258 116 265
rect 151 270 155 275
rect 151 268 152 270
rect 154 268 155 270
rect 95 245 97 247
rect 99 245 100 247
rect 95 240 100 245
rect 95 234 107 240
rect 151 247 155 268
rect 139 245 155 247
rect 139 243 141 245
rect 143 243 155 245
rect 139 242 155 243
rect 169 276 181 280
rect 169 274 171 276
rect 173 274 181 276
rect 245 278 269 279
rect 169 262 173 274
rect 245 276 247 278
rect 249 276 269 278
rect 245 275 269 276
rect 169 260 170 262
rect 172 260 173 262
rect 169 254 173 260
rect 193 271 198 272
rect 193 269 194 271
rect 196 269 198 271
rect 193 263 198 269
rect 169 252 174 254
rect 169 250 171 252
rect 173 250 174 252
rect 169 245 174 250
rect 169 243 171 245
rect 173 243 174 245
rect 184 262 198 263
rect 184 260 188 262
rect 190 260 198 262
rect 184 259 198 260
rect 217 271 230 272
rect 217 269 219 271
rect 221 269 230 271
rect 217 267 230 269
rect 217 266 227 267
rect 225 265 227 266
rect 229 265 230 267
rect 192 254 205 255
rect 192 252 198 254
rect 200 252 205 254
rect 192 251 205 252
rect 169 241 174 243
rect 201 247 205 251
rect 201 245 202 247
rect 204 245 205 247
rect 201 242 205 245
rect 209 254 214 256
rect 209 252 211 254
rect 213 252 214 254
rect 209 247 214 252
rect 225 258 230 265
rect 209 245 211 247
rect 213 245 214 247
rect 209 240 214 245
rect 209 234 221 240
rect 265 255 269 275
rect 287 263 292 272
rect 304 276 316 280
rect 304 274 312 276
rect 314 274 316 276
rect 287 262 301 263
rect 287 260 295 262
rect 297 260 301 262
rect 287 259 301 260
rect 265 253 266 255
rect 268 253 269 255
rect 265 247 269 253
rect 253 245 269 247
rect 253 243 255 245
rect 257 243 269 245
rect 253 242 269 243
rect 280 254 293 255
rect 280 252 285 254
rect 287 252 293 254
rect 280 251 293 252
rect 280 242 284 251
rect 312 270 316 274
rect 312 268 313 270
rect 315 268 316 270
rect 312 254 316 268
rect 311 252 316 254
rect 311 250 312 252
rect 314 250 316 252
rect 378 278 382 280
rect 377 276 382 278
rect 377 274 378 276
rect 380 274 382 276
rect 377 272 382 274
rect 329 270 342 271
rect 329 268 330 270
rect 332 268 342 270
rect 329 267 342 268
rect 336 262 342 267
rect 336 260 337 262
rect 339 260 342 262
rect 336 258 342 260
rect 362 257 366 264
rect 362 256 364 257
rect 354 255 364 256
rect 354 254 366 255
rect 354 252 355 254
rect 357 252 366 254
rect 354 250 366 252
rect 311 245 316 250
rect 311 243 312 245
rect 314 243 316 245
rect 311 241 316 243
rect 322 246 335 247
rect 322 244 332 246
rect 334 244 335 246
rect 322 243 335 244
rect 322 242 327 243
rect 378 262 382 272
rect 378 260 379 262
rect 381 260 382 262
rect 322 240 324 242
rect 326 240 327 242
rect 322 234 327 240
rect 378 239 382 260
rect 369 238 382 239
rect 369 236 378 238
rect 380 236 382 238
rect 369 235 382 236
rect 389 278 393 280
rect 389 276 394 278
rect 389 274 391 276
rect 393 274 394 276
rect 456 278 460 280
rect 389 272 394 274
rect 389 239 393 272
rect 429 270 442 271
rect 405 262 409 264
rect 405 260 406 262
rect 408 260 409 262
rect 405 257 409 260
rect 407 256 409 257
rect 407 255 417 256
rect 405 250 417 255
rect 429 268 437 270
rect 439 268 442 270
rect 429 267 442 268
rect 429 262 435 267
rect 429 260 432 262
rect 434 260 435 262
rect 429 258 435 260
rect 456 276 461 278
rect 456 274 458 276
rect 460 274 461 276
rect 564 278 588 279
rect 456 272 461 274
rect 456 270 460 272
rect 456 268 457 270
rect 459 268 460 270
rect 496 270 509 271
rect 436 243 449 247
rect 444 242 449 243
rect 389 238 402 239
rect 444 240 445 242
rect 447 240 449 242
rect 389 236 391 238
rect 393 236 402 238
rect 389 235 402 236
rect 444 234 449 240
rect 456 239 460 268
rect 472 257 476 264
rect 474 256 476 257
rect 474 255 484 256
rect 472 253 480 255
rect 482 253 484 255
rect 472 250 484 253
rect 496 268 505 270
rect 507 268 509 270
rect 496 267 509 268
rect 496 262 502 267
rect 496 260 499 262
rect 501 260 502 262
rect 496 258 502 260
rect 564 276 584 278
rect 586 276 588 278
rect 564 275 588 276
rect 522 271 527 273
rect 522 269 524 271
rect 526 269 527 271
rect 522 267 527 269
rect 522 254 526 267
rect 522 252 523 254
rect 525 252 526 254
rect 522 248 526 252
rect 554 263 558 272
rect 503 246 516 247
rect 503 244 504 246
rect 506 244 516 246
rect 503 243 516 244
rect 511 242 516 243
rect 456 238 469 239
rect 511 240 512 242
rect 514 240 516 242
rect 456 236 458 238
rect 460 236 469 238
rect 456 235 469 236
rect 511 234 516 240
rect 522 246 524 248
rect 522 241 526 246
rect 522 239 524 241
rect 537 262 558 263
rect 537 260 541 262
rect 543 260 558 262
rect 537 259 558 260
rect 564 270 568 275
rect 564 268 565 270
rect 567 268 568 270
rect 537 253 551 255
rect 553 253 558 255
rect 537 251 558 253
rect 554 242 558 251
rect 564 247 568 268
rect 603 267 616 272
rect 603 265 604 267
rect 606 266 616 267
rect 606 265 608 266
rect 564 245 580 247
rect 564 243 576 245
rect 578 243 580 245
rect 564 242 580 243
rect 603 258 608 265
rect 619 254 624 256
rect 619 252 620 254
rect 622 252 624 254
rect 522 235 535 239
rect 619 240 624 252
rect 522 234 526 235
rect 612 234 624 240
rect 2 228 632 229
rect 2 226 9 228
rect 11 226 58 228
rect 60 226 131 228
rect 133 226 172 228
rect 174 226 245 228
rect 247 226 311 228
rect 313 226 525 228
rect 527 226 586 228
rect 588 226 632 228
rect 2 216 632 226
rect 2 214 9 216
rect 11 214 58 216
rect 60 214 131 216
rect 133 214 172 216
rect 174 214 245 216
rect 247 214 311 216
rect 313 214 525 216
rect 527 214 586 216
rect 588 214 632 216
rect 2 213 632 214
rect 6 207 10 208
rect 6 203 19 207
rect 6 201 8 203
rect 6 196 10 201
rect 6 194 8 196
rect 6 175 10 194
rect 38 197 42 200
rect 55 199 60 201
rect 55 197 57 199
rect 59 197 60 199
rect 95 202 107 208
rect 38 193 60 197
rect 38 191 42 193
rect 21 189 42 191
rect 21 187 35 189
rect 37 187 42 189
rect 55 192 60 193
rect 55 190 57 192
rect 59 190 60 192
rect 55 188 60 190
rect 87 197 91 200
rect 87 195 88 197
rect 90 195 91 197
rect 6 173 11 175
rect 6 171 8 173
rect 10 171 11 173
rect 6 169 11 171
rect 21 182 42 183
rect 21 180 25 182
rect 27 180 39 182
rect 41 180 42 182
rect 21 179 42 180
rect 38 170 42 179
rect 55 168 59 188
rect 87 191 91 195
rect 78 190 91 191
rect 78 188 84 190
rect 86 188 91 190
rect 78 187 91 188
rect 95 197 100 202
rect 95 195 97 197
rect 99 195 100 197
rect 95 190 100 195
rect 95 188 97 190
rect 99 188 100 190
rect 95 186 100 188
rect 70 182 84 183
rect 70 180 74 182
rect 76 180 84 182
rect 70 179 84 180
rect 55 166 57 168
rect 59 166 67 168
rect 55 162 67 166
rect 79 173 84 179
rect 79 171 80 173
rect 82 171 84 173
rect 79 170 84 171
rect 111 177 116 184
rect 139 199 155 200
rect 139 197 141 199
rect 143 197 155 199
rect 139 195 155 197
rect 111 176 113 177
rect 103 175 113 176
rect 115 175 116 177
rect 103 173 116 175
rect 103 171 105 173
rect 107 171 116 173
rect 103 170 116 171
rect 151 174 155 195
rect 151 172 152 174
rect 154 172 155 174
rect 151 167 155 172
rect 131 166 155 167
rect 131 164 133 166
rect 135 164 155 166
rect 131 163 155 164
rect 169 199 174 201
rect 169 197 171 199
rect 173 197 174 199
rect 209 202 221 208
rect 169 192 174 197
rect 169 190 171 192
rect 173 190 174 192
rect 169 188 174 190
rect 201 197 205 200
rect 201 195 202 197
rect 204 195 205 197
rect 169 182 173 188
rect 169 180 170 182
rect 172 180 173 182
rect 169 168 173 180
rect 201 191 205 195
rect 192 190 205 191
rect 192 188 198 190
rect 200 188 205 190
rect 192 187 205 188
rect 209 197 214 202
rect 209 195 211 197
rect 213 195 214 197
rect 209 190 214 195
rect 209 188 211 190
rect 213 188 214 190
rect 209 186 214 188
rect 184 182 198 183
rect 184 180 188 182
rect 190 180 198 182
rect 184 179 198 180
rect 169 166 171 168
rect 173 166 181 168
rect 169 162 181 166
rect 193 173 198 179
rect 193 171 194 173
rect 196 171 198 173
rect 193 170 198 171
rect 225 177 230 184
rect 253 199 269 200
rect 253 197 255 199
rect 257 197 269 199
rect 253 195 269 197
rect 265 189 269 195
rect 265 187 266 189
rect 268 187 269 189
rect 280 191 284 200
rect 322 202 327 208
rect 369 206 382 207
rect 369 204 378 206
rect 380 204 382 206
rect 311 199 316 201
rect 280 190 293 191
rect 280 188 285 190
rect 287 188 293 190
rect 280 187 293 188
rect 225 176 227 177
rect 217 175 227 176
rect 229 175 230 177
rect 217 173 230 175
rect 217 171 219 173
rect 221 171 230 173
rect 217 170 230 171
rect 265 167 269 187
rect 287 182 301 183
rect 287 180 295 182
rect 297 180 301 182
rect 287 179 301 180
rect 311 197 312 199
rect 314 197 316 199
rect 311 192 316 197
rect 322 200 324 202
rect 326 200 327 202
rect 369 203 382 204
rect 322 199 327 200
rect 322 198 335 199
rect 322 196 332 198
rect 334 196 335 198
rect 322 195 335 196
rect 311 190 312 192
rect 314 190 316 192
rect 311 188 316 190
rect 287 170 292 179
rect 312 174 316 188
rect 312 172 313 174
rect 315 172 316 174
rect 312 168 316 172
rect 245 166 269 167
rect 245 164 247 166
rect 249 164 269 166
rect 245 163 269 164
rect 304 166 312 168
rect 314 166 316 168
rect 304 162 316 166
rect 336 182 342 184
rect 336 180 337 182
rect 339 180 342 182
rect 336 175 342 180
rect 329 174 342 175
rect 329 172 330 174
rect 332 172 342 174
rect 354 190 366 192
rect 354 188 355 190
rect 357 188 366 190
rect 354 187 366 188
rect 354 186 364 187
rect 362 185 364 186
rect 362 178 366 185
rect 378 182 382 203
rect 378 180 379 182
rect 381 180 382 182
rect 329 171 342 172
rect 378 170 382 180
rect 377 168 382 170
rect 377 166 378 168
rect 380 166 382 168
rect 377 164 382 166
rect 378 162 382 164
rect 389 206 402 207
rect 389 204 391 206
rect 393 204 402 206
rect 389 203 402 204
rect 389 170 393 203
rect 444 202 449 208
rect 444 200 445 202
rect 447 200 449 202
rect 444 199 449 200
rect 436 195 449 199
rect 456 206 469 207
rect 456 204 458 206
rect 460 204 469 206
rect 456 203 469 204
rect 405 187 417 192
rect 407 186 417 187
rect 407 185 409 186
rect 405 182 409 185
rect 405 180 406 182
rect 408 180 409 182
rect 405 178 409 180
rect 429 182 435 184
rect 429 180 432 182
rect 434 180 435 182
rect 429 175 435 180
rect 429 174 442 175
rect 429 172 437 174
rect 439 172 442 174
rect 429 171 442 172
rect 389 168 394 170
rect 389 166 391 168
rect 393 166 394 168
rect 389 164 394 166
rect 389 162 393 164
rect 456 174 460 203
rect 511 202 516 208
rect 511 200 512 202
rect 514 200 516 202
rect 511 199 516 200
rect 503 198 516 199
rect 503 196 504 198
rect 506 196 516 198
rect 503 195 516 196
rect 522 207 526 208
rect 522 203 535 207
rect 522 201 524 203
rect 522 196 526 201
rect 522 194 524 196
rect 472 189 484 192
rect 472 187 480 189
rect 482 187 484 189
rect 474 186 484 187
rect 474 185 476 186
rect 456 172 457 174
rect 459 172 460 174
rect 472 178 476 185
rect 456 170 460 172
rect 496 182 502 184
rect 496 180 499 182
rect 501 180 502 182
rect 496 175 502 180
rect 496 174 509 175
rect 496 172 505 174
rect 507 172 509 174
rect 496 171 509 172
rect 456 168 461 170
rect 456 166 458 168
rect 460 166 461 168
rect 456 164 461 166
rect 456 162 460 164
rect 522 190 526 194
rect 522 188 523 190
rect 525 188 526 190
rect 522 175 526 188
rect 554 191 558 200
rect 537 189 558 191
rect 537 187 551 189
rect 553 187 558 189
rect 564 199 580 200
rect 564 197 576 199
rect 578 197 580 199
rect 564 195 580 197
rect 522 173 527 175
rect 522 171 524 173
rect 526 171 527 173
rect 522 169 527 171
rect 537 182 558 183
rect 537 180 541 182
rect 543 180 558 182
rect 537 179 558 180
rect 554 170 558 179
rect 564 174 568 195
rect 612 202 624 208
rect 564 172 565 174
rect 567 172 568 174
rect 564 167 568 172
rect 603 177 608 184
rect 619 190 624 202
rect 619 188 620 190
rect 622 188 624 190
rect 619 186 624 188
rect 603 175 604 177
rect 606 176 608 177
rect 606 175 616 176
rect 603 170 616 175
rect 564 166 588 167
rect 564 164 584 166
rect 586 164 588 166
rect 564 163 588 164
rect 2 156 632 157
rect 2 154 9 156
rect 11 154 58 156
rect 60 154 68 156
rect 70 154 98 156
rect 100 154 151 156
rect 153 154 172 156
rect 174 154 182 156
rect 184 154 212 156
rect 214 154 265 156
rect 267 154 301 156
rect 303 154 311 156
rect 313 154 525 156
rect 527 154 566 156
rect 568 154 619 156
rect 621 154 632 156
rect 2 144 632 154
rect 2 142 9 144
rect 11 142 58 144
rect 60 142 68 144
rect 70 142 98 144
rect 100 142 151 144
rect 153 142 172 144
rect 174 142 182 144
rect 184 142 212 144
rect 214 142 265 144
rect 267 142 301 144
rect 303 142 311 144
rect 313 142 525 144
rect 527 142 566 144
rect 568 142 619 144
rect 621 142 632 144
rect 2 141 632 142
rect 55 132 67 136
rect 55 130 57 132
rect 59 130 67 132
rect 131 134 155 135
rect 6 127 11 129
rect 6 125 8 127
rect 10 125 11 127
rect 6 123 11 125
rect 6 104 10 123
rect 38 119 42 128
rect 6 102 8 104
rect 6 97 10 102
rect 6 95 8 97
rect 21 118 42 119
rect 21 116 25 118
rect 27 116 39 118
rect 41 116 42 118
rect 21 115 42 116
rect 21 109 35 111
rect 37 109 42 111
rect 21 107 42 109
rect 38 105 42 107
rect 55 110 59 130
rect 131 132 133 134
rect 135 132 155 134
rect 131 131 155 132
rect 79 127 84 128
rect 79 125 80 127
rect 82 125 84 127
rect 79 119 84 125
rect 55 108 60 110
rect 55 106 57 108
rect 59 106 60 108
rect 55 105 60 106
rect 38 101 60 105
rect 38 98 42 101
rect 55 99 57 101
rect 59 99 60 101
rect 70 118 84 119
rect 70 116 74 118
rect 76 116 84 118
rect 70 115 84 116
rect 103 127 116 128
rect 103 125 105 127
rect 107 125 116 127
rect 103 123 116 125
rect 103 122 113 123
rect 111 121 113 122
rect 115 121 116 123
rect 78 110 91 111
rect 78 108 84 110
rect 86 108 91 110
rect 78 107 91 108
rect 55 97 60 99
rect 6 91 19 95
rect 6 90 10 91
rect 87 103 91 107
rect 87 101 88 103
rect 90 101 91 103
rect 87 98 91 101
rect 95 110 100 112
rect 95 108 97 110
rect 99 108 100 110
rect 95 103 100 108
rect 111 114 116 121
rect 151 126 155 131
rect 151 124 152 126
rect 154 124 155 126
rect 95 101 97 103
rect 99 101 100 103
rect 95 96 100 101
rect 95 90 107 96
rect 151 103 155 124
rect 139 101 155 103
rect 139 99 141 101
rect 143 99 155 101
rect 139 98 155 99
rect 169 132 181 136
rect 169 130 171 132
rect 173 130 181 132
rect 245 134 269 135
rect 169 118 173 130
rect 245 132 247 134
rect 249 132 269 134
rect 245 131 269 132
rect 169 116 170 118
rect 172 116 173 118
rect 169 110 173 116
rect 193 127 198 128
rect 193 125 194 127
rect 196 125 198 127
rect 193 119 198 125
rect 169 108 174 110
rect 169 106 171 108
rect 173 106 174 108
rect 169 101 174 106
rect 169 99 171 101
rect 173 99 174 101
rect 184 118 198 119
rect 184 116 188 118
rect 190 116 198 118
rect 184 115 198 116
rect 217 127 230 128
rect 217 125 219 127
rect 221 125 230 127
rect 217 123 230 125
rect 217 122 227 123
rect 225 121 227 122
rect 229 121 230 123
rect 192 110 205 111
rect 192 108 198 110
rect 200 108 205 110
rect 192 107 205 108
rect 169 97 174 99
rect 201 103 205 107
rect 201 101 202 103
rect 204 101 205 103
rect 201 98 205 101
rect 209 110 214 112
rect 209 108 211 110
rect 213 108 214 110
rect 209 103 214 108
rect 225 114 230 121
rect 209 101 211 103
rect 213 101 214 103
rect 209 96 214 101
rect 209 90 221 96
rect 265 111 269 131
rect 287 119 292 128
rect 304 132 316 136
rect 304 130 312 132
rect 314 130 316 132
rect 287 118 301 119
rect 287 116 295 118
rect 297 116 301 118
rect 287 115 301 116
rect 265 109 266 111
rect 268 109 269 111
rect 265 103 269 109
rect 253 101 269 103
rect 253 99 255 101
rect 257 99 269 101
rect 253 98 269 99
rect 280 110 293 111
rect 280 108 285 110
rect 287 108 293 110
rect 280 107 293 108
rect 280 98 284 107
rect 312 126 316 130
rect 312 124 313 126
rect 315 124 316 126
rect 312 110 316 124
rect 311 108 316 110
rect 311 106 312 108
rect 314 106 316 108
rect 378 134 382 136
rect 377 132 382 134
rect 377 130 378 132
rect 380 130 382 132
rect 377 128 382 130
rect 329 126 342 127
rect 329 124 330 126
rect 332 124 342 126
rect 329 123 342 124
rect 336 118 342 123
rect 336 116 337 118
rect 339 116 342 118
rect 336 114 342 116
rect 362 113 366 120
rect 362 112 364 113
rect 354 111 364 112
rect 354 110 366 111
rect 354 108 355 110
rect 357 108 366 110
rect 354 106 366 108
rect 311 101 316 106
rect 311 99 312 101
rect 314 99 316 101
rect 311 97 316 99
rect 322 102 335 103
rect 322 100 332 102
rect 334 100 335 102
rect 322 99 335 100
rect 322 98 327 99
rect 378 118 382 128
rect 378 116 379 118
rect 381 116 382 118
rect 322 96 324 98
rect 326 96 327 98
rect 322 90 327 96
rect 378 95 382 116
rect 369 94 382 95
rect 369 92 378 94
rect 380 92 382 94
rect 369 91 382 92
rect 389 134 393 136
rect 389 132 394 134
rect 389 130 391 132
rect 393 130 394 132
rect 456 134 460 136
rect 389 128 394 130
rect 389 95 393 128
rect 429 126 442 127
rect 405 118 409 120
rect 405 116 406 118
rect 408 116 409 118
rect 405 113 409 116
rect 407 112 409 113
rect 407 111 417 112
rect 405 106 417 111
rect 429 124 437 126
rect 439 124 442 126
rect 429 123 442 124
rect 429 118 435 123
rect 429 116 432 118
rect 434 116 435 118
rect 429 114 435 116
rect 456 132 461 134
rect 456 130 458 132
rect 460 130 461 132
rect 564 134 588 135
rect 456 128 461 130
rect 456 126 460 128
rect 456 124 457 126
rect 459 124 460 126
rect 496 126 509 127
rect 436 99 449 103
rect 444 98 449 99
rect 389 94 402 95
rect 444 96 445 98
rect 447 96 449 98
rect 389 92 391 94
rect 393 92 402 94
rect 389 91 402 92
rect 444 90 449 96
rect 456 95 460 124
rect 472 113 476 120
rect 474 112 476 113
rect 474 111 484 112
rect 472 109 480 111
rect 482 109 484 111
rect 472 106 484 109
rect 496 124 505 126
rect 507 124 509 126
rect 496 123 509 124
rect 496 118 502 123
rect 496 116 499 118
rect 501 116 502 118
rect 496 114 502 116
rect 564 132 584 134
rect 586 132 588 134
rect 564 131 588 132
rect 522 127 527 129
rect 522 125 524 127
rect 526 125 527 127
rect 522 123 527 125
rect 522 110 526 123
rect 522 108 523 110
rect 525 108 526 110
rect 522 104 526 108
rect 554 119 558 128
rect 503 102 516 103
rect 503 100 504 102
rect 506 100 516 102
rect 503 99 516 100
rect 511 98 516 99
rect 456 94 469 95
rect 511 96 512 98
rect 514 96 516 98
rect 456 92 458 94
rect 460 92 469 94
rect 456 91 469 92
rect 511 90 516 96
rect 522 102 524 104
rect 522 97 526 102
rect 522 95 524 97
rect 537 118 558 119
rect 537 116 541 118
rect 543 116 558 118
rect 537 115 558 116
rect 564 126 568 131
rect 564 124 565 126
rect 567 124 568 126
rect 537 109 551 111
rect 553 109 558 111
rect 537 107 558 109
rect 554 98 558 107
rect 564 103 568 124
rect 603 123 616 128
rect 603 121 604 123
rect 606 122 616 123
rect 606 121 608 122
rect 564 101 580 103
rect 564 99 576 101
rect 578 99 580 101
rect 564 98 580 99
rect 603 114 608 121
rect 619 110 624 112
rect 619 108 620 110
rect 622 108 624 110
rect 522 91 535 95
rect 619 96 624 108
rect 522 90 526 91
rect 612 90 624 96
rect 2 84 632 85
rect 2 82 9 84
rect 11 82 58 84
rect 60 82 131 84
rect 133 82 172 84
rect 174 82 245 84
rect 247 82 311 84
rect 313 82 525 84
rect 527 82 586 84
rect 588 82 632 84
rect 2 72 632 82
rect 2 70 9 72
rect 11 70 58 72
rect 60 70 131 72
rect 133 70 172 72
rect 174 70 245 72
rect 247 70 311 72
rect 313 70 525 72
rect 527 70 586 72
rect 588 70 632 72
rect 2 69 632 70
rect 6 63 10 64
rect 6 59 19 63
rect 6 57 8 59
rect 6 52 10 57
rect 6 50 8 52
rect 6 31 10 50
rect 38 53 42 56
rect 55 55 60 57
rect 55 53 57 55
rect 59 53 60 55
rect 95 58 107 64
rect 38 49 60 53
rect 38 47 42 49
rect 21 45 42 47
rect 21 43 35 45
rect 37 43 42 45
rect 55 48 60 49
rect 55 46 57 48
rect 59 46 60 48
rect 55 44 60 46
rect 87 53 91 56
rect 87 51 88 53
rect 90 51 91 53
rect 6 29 11 31
rect 6 27 8 29
rect 10 27 11 29
rect 6 25 11 27
rect 21 38 42 39
rect 21 36 25 38
rect 27 36 39 38
rect 41 36 42 38
rect 21 35 42 36
rect 38 26 42 35
rect 55 24 59 44
rect 87 47 91 51
rect 78 46 91 47
rect 78 44 84 46
rect 86 44 91 46
rect 78 43 91 44
rect 95 53 100 58
rect 95 51 97 53
rect 99 51 100 53
rect 95 46 100 51
rect 95 44 97 46
rect 99 44 100 46
rect 95 42 100 44
rect 70 38 84 39
rect 70 36 74 38
rect 76 36 84 38
rect 70 35 84 36
rect 55 22 57 24
rect 59 22 67 24
rect 55 18 67 22
rect 79 29 84 35
rect 79 27 80 29
rect 82 27 84 29
rect 79 26 84 27
rect 111 33 116 40
rect 139 55 155 56
rect 139 53 141 55
rect 143 53 155 55
rect 139 51 155 53
rect 111 32 113 33
rect 103 31 113 32
rect 115 31 116 33
rect 103 29 116 31
rect 103 27 105 29
rect 107 27 116 29
rect 103 26 116 27
rect 151 30 155 51
rect 151 28 152 30
rect 154 28 155 30
rect 151 23 155 28
rect 131 22 155 23
rect 131 20 133 22
rect 135 20 155 22
rect 131 19 155 20
rect 169 55 174 57
rect 169 53 171 55
rect 173 53 174 55
rect 209 58 221 64
rect 169 48 174 53
rect 169 46 171 48
rect 173 46 174 48
rect 169 44 174 46
rect 201 53 205 56
rect 201 51 202 53
rect 204 51 205 53
rect 169 38 173 44
rect 169 36 170 38
rect 172 36 173 38
rect 169 24 173 36
rect 201 47 205 51
rect 192 46 205 47
rect 192 44 198 46
rect 200 44 205 46
rect 192 43 205 44
rect 209 53 214 58
rect 209 51 211 53
rect 213 51 214 53
rect 209 46 214 51
rect 209 44 211 46
rect 213 44 214 46
rect 209 42 214 44
rect 184 38 198 39
rect 184 36 188 38
rect 190 36 198 38
rect 184 35 198 36
rect 169 22 171 24
rect 173 22 181 24
rect 169 18 181 22
rect 193 29 198 35
rect 193 27 194 29
rect 196 27 198 29
rect 193 26 198 27
rect 225 33 230 40
rect 253 55 269 56
rect 253 53 255 55
rect 257 53 269 55
rect 253 51 269 53
rect 265 45 269 51
rect 265 43 266 45
rect 268 43 269 45
rect 280 47 284 56
rect 322 58 327 64
rect 369 62 382 63
rect 369 60 378 62
rect 380 60 382 62
rect 311 55 316 57
rect 280 46 293 47
rect 280 44 285 46
rect 287 44 293 46
rect 280 43 293 44
rect 225 32 227 33
rect 217 31 227 32
rect 229 31 230 33
rect 217 29 230 31
rect 217 27 219 29
rect 221 27 230 29
rect 217 26 230 27
rect 265 23 269 43
rect 287 38 301 39
rect 287 36 295 38
rect 297 36 301 38
rect 287 35 301 36
rect 311 53 312 55
rect 314 53 316 55
rect 311 48 316 53
rect 322 56 324 58
rect 326 56 327 58
rect 369 59 382 60
rect 322 55 327 56
rect 322 54 335 55
rect 322 52 332 54
rect 334 52 335 54
rect 322 51 335 52
rect 311 46 312 48
rect 314 46 316 48
rect 311 44 316 46
rect 287 26 292 35
rect 312 30 316 44
rect 312 28 313 30
rect 315 28 316 30
rect 312 24 316 28
rect 245 22 269 23
rect 245 20 247 22
rect 249 20 269 22
rect 245 19 269 20
rect 304 22 312 24
rect 314 22 316 24
rect 304 18 316 22
rect 336 38 342 40
rect 336 36 337 38
rect 339 36 342 38
rect 336 31 342 36
rect 329 30 342 31
rect 329 28 330 30
rect 332 28 342 30
rect 354 46 366 48
rect 354 44 355 46
rect 357 44 366 46
rect 354 43 366 44
rect 354 42 364 43
rect 362 41 364 42
rect 362 34 366 41
rect 378 38 382 59
rect 378 36 379 38
rect 381 36 382 38
rect 329 27 342 28
rect 378 26 382 36
rect 377 24 382 26
rect 377 22 378 24
rect 380 22 382 24
rect 377 20 382 22
rect 378 18 382 20
rect 389 62 402 63
rect 389 60 391 62
rect 393 60 402 62
rect 389 59 402 60
rect 389 26 393 59
rect 444 58 449 64
rect 444 56 445 58
rect 447 56 449 58
rect 444 55 449 56
rect 436 51 449 55
rect 456 62 469 63
rect 456 60 458 62
rect 460 60 469 62
rect 456 59 469 60
rect 405 43 417 48
rect 407 42 417 43
rect 407 41 409 42
rect 405 38 409 41
rect 405 36 406 38
rect 408 36 409 38
rect 405 34 409 36
rect 429 38 435 40
rect 429 36 432 38
rect 434 36 435 38
rect 429 31 435 36
rect 429 30 442 31
rect 429 28 437 30
rect 439 28 442 30
rect 429 27 442 28
rect 389 24 394 26
rect 389 22 391 24
rect 393 22 394 24
rect 389 20 394 22
rect 389 18 393 20
rect 456 30 460 59
rect 511 58 516 64
rect 511 56 512 58
rect 514 56 516 58
rect 511 55 516 56
rect 503 54 516 55
rect 503 52 504 54
rect 506 52 516 54
rect 503 51 516 52
rect 522 63 526 64
rect 522 59 535 63
rect 522 57 524 59
rect 522 52 526 57
rect 522 50 524 52
rect 472 45 484 48
rect 472 43 480 45
rect 482 43 484 45
rect 474 42 484 43
rect 474 41 476 42
rect 456 28 457 30
rect 459 28 460 30
rect 472 34 476 41
rect 456 26 460 28
rect 496 38 502 40
rect 496 36 499 38
rect 501 36 502 38
rect 496 31 502 36
rect 496 30 509 31
rect 496 28 505 30
rect 507 28 509 30
rect 496 27 509 28
rect 456 24 461 26
rect 456 22 458 24
rect 460 22 461 24
rect 456 20 461 22
rect 456 18 460 20
rect 522 46 526 50
rect 522 44 523 46
rect 525 44 526 46
rect 522 31 526 44
rect 554 47 558 56
rect 537 45 558 47
rect 537 43 551 45
rect 553 43 558 45
rect 564 55 580 56
rect 564 53 576 55
rect 578 53 580 55
rect 564 51 580 53
rect 522 29 527 31
rect 522 27 524 29
rect 526 27 527 29
rect 522 25 527 27
rect 537 38 558 39
rect 537 36 541 38
rect 543 36 558 38
rect 537 35 558 36
rect 554 26 558 35
rect 564 30 568 51
rect 612 58 624 64
rect 564 28 565 30
rect 567 28 568 30
rect 564 23 568 28
rect 603 33 608 40
rect 619 46 624 58
rect 619 44 620 46
rect 622 44 624 46
rect 619 42 624 44
rect 603 31 604 33
rect 606 32 608 33
rect 606 31 616 32
rect 603 26 616 31
rect 564 22 588 23
rect 564 20 584 22
rect 586 20 588 22
rect 564 19 588 20
rect 2 12 632 13
rect 2 10 9 12
rect 11 10 58 12
rect 60 10 68 12
rect 70 10 98 12
rect 100 10 151 12
rect 153 10 172 12
rect 174 10 182 12
rect 184 10 212 12
rect 214 10 265 12
rect 267 10 301 12
rect 303 10 311 12
rect 313 10 525 12
rect 527 10 566 12
rect 568 10 619 12
rect 621 10 632 12
rect 2 5 632 10
<< alu2 >>
rect 79 559 111 560
rect 79 557 80 559
rect 82 557 105 559
rect 107 557 111 559
rect 79 555 111 557
rect 151 559 225 560
rect 151 558 194 559
rect 151 556 152 558
rect 154 557 194 558
rect 196 557 219 559
rect 221 557 225 559
rect 154 556 225 557
rect 151 555 225 556
rect 312 558 333 559
rect 312 556 313 558
rect 315 556 330 558
rect 332 556 333 558
rect 312 555 333 556
rect 436 558 460 559
rect 436 556 437 558
rect 439 556 457 558
rect 459 556 460 558
rect 436 555 460 556
rect 504 558 568 559
rect 504 556 505 558
rect 507 556 565 558
rect 567 556 568 558
rect 504 555 568 556
rect 38 550 173 551
rect 38 548 39 550
rect 41 548 170 550
rect 172 548 173 550
rect 38 547 173 548
rect 378 550 409 551
rect 378 548 379 550
rect 381 548 406 550
rect 408 548 409 550
rect 378 547 409 548
rect 265 543 359 544
rect 265 541 266 543
rect 268 542 359 543
rect 268 541 355 542
rect 265 540 355 541
rect 357 540 359 542
rect 265 539 359 540
rect 479 543 526 544
rect 479 541 480 543
rect 482 542 526 543
rect 482 541 523 542
rect 479 540 523 541
rect 525 540 526 542
rect 479 539 526 540
rect 87 535 100 536
rect 87 533 88 535
rect 90 533 97 535
rect 99 533 100 535
rect 87 532 100 533
rect 201 535 214 536
rect 201 533 202 535
rect 204 533 211 535
rect 213 533 214 535
rect 201 532 214 533
rect 331 534 508 535
rect 331 532 332 534
rect 334 532 504 534
rect 506 532 508 534
rect 331 531 508 532
rect 331 486 508 487
rect 87 485 100 486
rect 87 483 88 485
rect 90 483 97 485
rect 99 483 100 485
rect 87 482 100 483
rect 201 485 214 486
rect 201 483 202 485
rect 204 483 211 485
rect 213 483 214 485
rect 331 484 332 486
rect 334 484 504 486
rect 506 484 508 486
rect 331 483 508 484
rect 201 482 214 483
rect 265 478 359 479
rect 265 477 355 478
rect 265 475 266 477
rect 268 476 355 477
rect 357 476 359 478
rect 268 475 359 476
rect 265 474 359 475
rect 479 478 526 479
rect 479 477 523 478
rect 479 475 480 477
rect 482 476 523 477
rect 525 476 526 478
rect 482 475 526 476
rect 479 474 526 475
rect 38 470 173 471
rect 38 468 39 470
rect 41 468 170 470
rect 172 468 173 470
rect 38 467 173 468
rect 378 470 409 471
rect 378 468 379 470
rect 381 468 406 470
rect 408 468 409 470
rect 378 467 409 468
rect 79 461 111 463
rect 79 459 80 461
rect 82 459 105 461
rect 107 459 111 461
rect 79 458 111 459
rect 151 462 225 463
rect 151 460 152 462
rect 154 461 225 462
rect 154 460 194 461
rect 151 459 194 460
rect 196 459 219 461
rect 221 459 225 461
rect 312 462 333 463
rect 312 460 313 462
rect 315 460 330 462
rect 332 460 333 462
rect 312 459 333 460
rect 436 462 460 463
rect 436 460 437 462
rect 439 460 457 462
rect 459 460 460 462
rect 436 459 460 460
rect 504 462 568 463
rect 504 460 505 462
rect 507 460 565 462
rect 567 460 568 462
rect 504 459 568 460
rect 151 458 225 459
rect 79 415 111 416
rect 79 413 80 415
rect 82 413 105 415
rect 107 413 111 415
rect 79 411 111 413
rect 151 415 225 416
rect 151 414 194 415
rect 151 412 152 414
rect 154 413 194 414
rect 196 413 219 415
rect 221 413 225 415
rect 154 412 225 413
rect 151 411 225 412
rect 312 414 333 415
rect 312 412 313 414
rect 315 412 330 414
rect 332 412 333 414
rect 312 411 333 412
rect 436 414 460 415
rect 436 412 437 414
rect 439 412 457 414
rect 459 412 460 414
rect 436 411 460 412
rect 504 414 568 415
rect 504 412 505 414
rect 507 412 565 414
rect 567 412 568 414
rect 504 411 568 412
rect 38 406 173 407
rect 38 404 39 406
rect 41 404 170 406
rect 172 404 173 406
rect 38 403 173 404
rect 378 406 409 407
rect 378 404 379 406
rect 381 404 406 406
rect 408 404 409 406
rect 378 403 409 404
rect 265 399 359 400
rect 265 397 266 399
rect 268 398 359 399
rect 268 397 355 398
rect 265 396 355 397
rect 357 396 359 398
rect 265 395 359 396
rect 479 399 526 400
rect 479 397 480 399
rect 482 398 526 399
rect 482 397 523 398
rect 479 396 523 397
rect 525 396 526 398
rect 479 395 526 396
rect 87 391 100 392
rect 87 389 88 391
rect 90 389 97 391
rect 99 389 100 391
rect 87 388 100 389
rect 201 391 214 392
rect 201 389 202 391
rect 204 389 211 391
rect 213 389 214 391
rect 201 388 214 389
rect 331 390 508 391
rect 331 388 332 390
rect 334 388 504 390
rect 506 388 508 390
rect 331 387 508 388
rect 331 342 508 343
rect 87 341 100 342
rect 87 339 88 341
rect 90 339 97 341
rect 99 339 100 341
rect 87 338 100 339
rect 201 341 214 342
rect 201 339 202 341
rect 204 339 211 341
rect 213 339 214 341
rect 331 340 332 342
rect 334 340 504 342
rect 506 340 508 342
rect 331 339 508 340
rect 201 338 214 339
rect 265 334 359 335
rect 265 333 355 334
rect 265 331 266 333
rect 268 332 355 333
rect 357 332 359 334
rect 268 331 359 332
rect 265 330 359 331
rect 479 334 526 335
rect 479 333 523 334
rect 479 331 480 333
rect 482 332 523 333
rect 525 332 526 334
rect 482 331 526 332
rect 479 330 526 331
rect 38 326 173 327
rect 38 324 39 326
rect 41 324 170 326
rect 172 324 173 326
rect 38 323 173 324
rect 378 326 409 327
rect 378 324 379 326
rect 381 324 406 326
rect 408 324 409 326
rect 378 323 409 324
rect 79 317 111 319
rect 79 315 80 317
rect 82 315 105 317
rect 107 315 111 317
rect 79 314 111 315
rect 151 318 225 319
rect 151 316 152 318
rect 154 317 225 318
rect 154 316 194 317
rect 151 315 194 316
rect 196 315 219 317
rect 221 315 225 317
rect 312 318 333 319
rect 312 316 313 318
rect 315 316 330 318
rect 332 316 333 318
rect 312 315 333 316
rect 436 318 460 319
rect 436 316 437 318
rect 439 316 457 318
rect 459 316 460 318
rect 436 315 460 316
rect 504 318 568 319
rect 504 316 505 318
rect 507 316 565 318
rect 567 316 568 318
rect 504 315 568 316
rect 151 314 225 315
rect 79 271 111 272
rect 79 269 80 271
rect 82 269 105 271
rect 107 269 111 271
rect 79 267 111 269
rect 151 271 225 272
rect 151 270 194 271
rect 151 268 152 270
rect 154 269 194 270
rect 196 269 219 271
rect 221 269 225 271
rect 154 268 225 269
rect 151 267 225 268
rect 312 270 333 271
rect 312 268 313 270
rect 315 268 330 270
rect 332 268 333 270
rect 312 267 333 268
rect 436 270 460 271
rect 436 268 437 270
rect 439 268 457 270
rect 459 268 460 270
rect 436 267 460 268
rect 504 270 568 271
rect 504 268 505 270
rect 507 268 565 270
rect 567 268 568 270
rect 504 267 568 268
rect 38 262 173 263
rect 38 260 39 262
rect 41 260 170 262
rect 172 260 173 262
rect 38 259 173 260
rect 378 262 409 263
rect 378 260 379 262
rect 381 260 406 262
rect 408 260 409 262
rect 378 259 409 260
rect 265 255 359 256
rect 265 253 266 255
rect 268 254 359 255
rect 268 253 355 254
rect 265 252 355 253
rect 357 252 359 254
rect 265 251 359 252
rect 479 255 526 256
rect 479 253 480 255
rect 482 254 526 255
rect 482 253 523 254
rect 479 252 523 253
rect 525 252 526 254
rect 479 251 526 252
rect 87 247 100 248
rect 87 245 88 247
rect 90 245 97 247
rect 99 245 100 247
rect 87 244 100 245
rect 201 247 214 248
rect 201 245 202 247
rect 204 245 211 247
rect 213 245 214 247
rect 201 244 214 245
rect 331 246 508 247
rect 331 244 332 246
rect 334 244 504 246
rect 506 244 508 246
rect 331 243 508 244
rect 331 198 508 199
rect 87 197 100 198
rect 87 195 88 197
rect 90 195 97 197
rect 99 195 100 197
rect 87 194 100 195
rect 201 197 214 198
rect 201 195 202 197
rect 204 195 211 197
rect 213 195 214 197
rect 331 196 332 198
rect 334 196 504 198
rect 506 196 508 198
rect 331 195 508 196
rect 201 194 214 195
rect 265 190 359 191
rect 265 189 355 190
rect 265 187 266 189
rect 268 188 355 189
rect 357 188 359 190
rect 268 187 359 188
rect 265 186 359 187
rect 479 190 526 191
rect 479 189 523 190
rect 479 187 480 189
rect 482 188 523 189
rect 525 188 526 190
rect 482 187 526 188
rect 479 186 526 187
rect 38 182 173 183
rect 38 180 39 182
rect 41 180 170 182
rect 172 180 173 182
rect 38 179 173 180
rect 378 182 409 183
rect 378 180 379 182
rect 381 180 406 182
rect 408 180 409 182
rect 378 179 409 180
rect 79 173 111 175
rect 79 171 80 173
rect 82 171 105 173
rect 107 171 111 173
rect 79 170 111 171
rect 151 174 225 175
rect 151 172 152 174
rect 154 173 225 174
rect 154 172 194 173
rect 151 171 194 172
rect 196 171 219 173
rect 221 171 225 173
rect 312 174 333 175
rect 312 172 313 174
rect 315 172 330 174
rect 332 172 333 174
rect 312 171 333 172
rect 436 174 460 175
rect 436 172 437 174
rect 439 172 457 174
rect 459 172 460 174
rect 436 171 460 172
rect 504 174 568 175
rect 504 172 505 174
rect 507 172 565 174
rect 567 172 568 174
rect 504 171 568 172
rect 151 170 225 171
rect 79 127 111 128
rect 79 125 80 127
rect 82 125 105 127
rect 107 125 111 127
rect 79 123 111 125
rect 151 127 225 128
rect 151 126 194 127
rect 151 124 152 126
rect 154 125 194 126
rect 196 125 219 127
rect 221 125 225 127
rect 154 124 225 125
rect 151 123 225 124
rect 312 126 333 127
rect 312 124 313 126
rect 315 124 330 126
rect 332 124 333 126
rect 312 123 333 124
rect 436 126 460 127
rect 436 124 437 126
rect 439 124 457 126
rect 459 124 460 126
rect 436 123 460 124
rect 504 126 568 127
rect 504 124 505 126
rect 507 124 565 126
rect 567 124 568 126
rect 504 123 568 124
rect 38 118 173 119
rect 38 116 39 118
rect 41 116 170 118
rect 172 116 173 118
rect 38 115 173 116
rect 378 118 409 119
rect 378 116 379 118
rect 381 116 406 118
rect 408 116 409 118
rect 378 115 409 116
rect 265 111 359 112
rect 265 109 266 111
rect 268 110 359 111
rect 268 109 355 110
rect 265 108 355 109
rect 357 108 359 110
rect 265 107 359 108
rect 479 111 526 112
rect 479 109 480 111
rect 482 110 526 111
rect 482 109 523 110
rect 479 108 523 109
rect 525 108 526 110
rect 479 107 526 108
rect 87 103 100 104
rect 87 101 88 103
rect 90 101 97 103
rect 99 101 100 103
rect 87 100 100 101
rect 201 103 214 104
rect 201 101 202 103
rect 204 101 211 103
rect 213 101 214 103
rect 201 100 214 101
rect 331 102 508 103
rect 331 100 332 102
rect 334 100 504 102
rect 506 100 508 102
rect 331 99 508 100
rect 331 54 508 55
rect 87 53 100 54
rect 87 51 88 53
rect 90 51 97 53
rect 99 51 100 53
rect 87 50 100 51
rect 201 53 214 54
rect 201 51 202 53
rect 204 51 211 53
rect 213 51 214 53
rect 331 52 332 54
rect 334 52 504 54
rect 506 52 508 54
rect 331 51 508 52
rect 201 50 214 51
rect 265 46 359 47
rect 265 45 355 46
rect 265 43 266 45
rect 268 44 355 45
rect 357 44 359 46
rect 268 43 359 44
rect 265 42 359 43
rect 479 46 526 47
rect 479 45 523 46
rect 479 43 480 45
rect 482 44 523 45
rect 525 44 526 46
rect 482 43 526 44
rect 479 42 526 43
rect 38 38 173 39
rect 38 36 39 38
rect 41 36 170 38
rect 172 36 173 38
rect 38 35 173 36
rect 378 38 409 39
rect 378 36 379 38
rect 381 36 406 38
rect 408 36 409 38
rect 378 35 409 36
rect 79 29 111 31
rect 79 27 80 29
rect 82 27 105 29
rect 107 27 111 29
rect 79 26 111 27
rect 151 30 225 31
rect 151 28 152 30
rect 154 29 225 30
rect 154 28 194 29
rect 151 27 194 28
rect 196 27 219 29
rect 221 27 225 29
rect 312 30 333 31
rect 312 28 313 30
rect 315 28 330 30
rect 332 28 333 30
rect 312 27 333 28
rect 436 30 460 31
rect 436 28 437 30
rect 439 28 457 30
rect 459 28 460 30
rect 436 27 460 28
rect 504 30 568 31
rect 504 28 505 30
rect 507 28 565 30
rect 567 28 568 30
rect 504 27 568 28
rect 151 26 225 27
<< ptie >>
rect 7 576 13 578
rect 7 574 9 576
rect 11 574 13 576
rect 56 576 62 578
rect 56 574 58 576
rect 60 574 62 576
rect 7 572 13 574
rect 56 572 62 574
rect 96 576 102 578
rect 96 574 98 576
rect 100 574 102 576
rect 96 572 102 574
rect 170 576 176 578
rect 170 574 172 576
rect 174 574 176 576
rect 170 572 176 574
rect 210 576 216 578
rect 210 574 212 576
rect 214 574 216 576
rect 210 572 216 574
rect 309 576 315 578
rect 309 574 311 576
rect 313 574 315 576
rect 309 572 315 574
rect 523 576 529 578
rect 523 574 525 576
rect 527 574 529 576
rect 523 572 529 574
rect 617 576 623 578
rect 617 574 619 576
rect 621 574 623 576
rect 617 572 623 574
rect 7 444 13 446
rect 56 444 62 446
rect 7 442 9 444
rect 11 442 13 444
rect 7 440 13 442
rect 56 442 58 444
rect 60 442 62 444
rect 56 440 62 442
rect 96 444 102 446
rect 96 442 98 444
rect 100 442 102 444
rect 96 440 102 442
rect 170 444 176 446
rect 170 442 172 444
rect 174 442 176 444
rect 170 440 176 442
rect 210 444 216 446
rect 210 442 212 444
rect 214 442 216 444
rect 210 440 216 442
rect 309 444 315 446
rect 309 442 311 444
rect 313 442 315 444
rect 309 440 315 442
rect 523 444 529 446
rect 523 442 525 444
rect 527 442 529 444
rect 523 440 529 442
rect 617 444 623 446
rect 617 442 619 444
rect 621 442 623 444
rect 617 440 623 442
rect 7 432 13 434
rect 7 430 9 432
rect 11 430 13 432
rect 56 432 62 434
rect 56 430 58 432
rect 60 430 62 432
rect 7 428 13 430
rect 56 428 62 430
rect 96 432 102 434
rect 96 430 98 432
rect 100 430 102 432
rect 96 428 102 430
rect 170 432 176 434
rect 170 430 172 432
rect 174 430 176 432
rect 170 428 176 430
rect 210 432 216 434
rect 210 430 212 432
rect 214 430 216 432
rect 210 428 216 430
rect 309 432 315 434
rect 309 430 311 432
rect 313 430 315 432
rect 309 428 315 430
rect 523 432 529 434
rect 523 430 525 432
rect 527 430 529 432
rect 523 428 529 430
rect 617 432 623 434
rect 617 430 619 432
rect 621 430 623 432
rect 617 428 623 430
rect 7 300 13 302
rect 56 300 62 302
rect 7 298 9 300
rect 11 298 13 300
rect 7 296 13 298
rect 56 298 58 300
rect 60 298 62 300
rect 56 296 62 298
rect 96 300 102 302
rect 96 298 98 300
rect 100 298 102 300
rect 96 296 102 298
rect 170 300 176 302
rect 170 298 172 300
rect 174 298 176 300
rect 170 296 176 298
rect 210 300 216 302
rect 210 298 212 300
rect 214 298 216 300
rect 210 296 216 298
rect 309 300 315 302
rect 309 298 311 300
rect 313 298 315 300
rect 309 296 315 298
rect 523 300 529 302
rect 523 298 525 300
rect 527 298 529 300
rect 523 296 529 298
rect 617 300 623 302
rect 617 298 619 300
rect 621 298 623 300
rect 617 296 623 298
rect 7 288 13 290
rect 7 286 9 288
rect 11 286 13 288
rect 56 288 62 290
rect 56 286 58 288
rect 60 286 62 288
rect 7 284 13 286
rect 56 284 62 286
rect 96 288 102 290
rect 96 286 98 288
rect 100 286 102 288
rect 96 284 102 286
rect 170 288 176 290
rect 170 286 172 288
rect 174 286 176 288
rect 170 284 176 286
rect 210 288 216 290
rect 210 286 212 288
rect 214 286 216 288
rect 210 284 216 286
rect 309 288 315 290
rect 309 286 311 288
rect 313 286 315 288
rect 309 284 315 286
rect 523 288 529 290
rect 523 286 525 288
rect 527 286 529 288
rect 523 284 529 286
rect 617 288 623 290
rect 617 286 619 288
rect 621 286 623 288
rect 617 284 623 286
rect 7 156 13 158
rect 56 156 62 158
rect 7 154 9 156
rect 11 154 13 156
rect 7 152 13 154
rect 56 154 58 156
rect 60 154 62 156
rect 56 152 62 154
rect 96 156 102 158
rect 96 154 98 156
rect 100 154 102 156
rect 96 152 102 154
rect 170 156 176 158
rect 170 154 172 156
rect 174 154 176 156
rect 170 152 176 154
rect 210 156 216 158
rect 210 154 212 156
rect 214 154 216 156
rect 210 152 216 154
rect 309 156 315 158
rect 309 154 311 156
rect 313 154 315 156
rect 309 152 315 154
rect 523 156 529 158
rect 523 154 525 156
rect 527 154 529 156
rect 523 152 529 154
rect 617 156 623 158
rect 617 154 619 156
rect 621 154 623 156
rect 617 152 623 154
rect 7 144 13 146
rect 7 142 9 144
rect 11 142 13 144
rect 56 144 62 146
rect 56 142 58 144
rect 60 142 62 144
rect 7 140 13 142
rect 56 140 62 142
rect 96 144 102 146
rect 96 142 98 144
rect 100 142 102 144
rect 96 140 102 142
rect 170 144 176 146
rect 170 142 172 144
rect 174 142 176 144
rect 170 140 176 142
rect 210 144 216 146
rect 210 142 212 144
rect 214 142 216 144
rect 210 140 216 142
rect 309 144 315 146
rect 309 142 311 144
rect 313 142 315 144
rect 309 140 315 142
rect 523 144 529 146
rect 523 142 525 144
rect 527 142 529 144
rect 523 140 529 142
rect 617 144 623 146
rect 617 142 619 144
rect 621 142 623 144
rect 617 140 623 142
rect 7 12 13 14
rect 56 12 62 14
rect 7 10 9 12
rect 11 10 13 12
rect 7 8 13 10
rect 56 10 58 12
rect 60 10 62 12
rect 56 8 62 10
rect 96 12 102 14
rect 96 10 98 12
rect 100 10 102 12
rect 96 8 102 10
rect 170 12 176 14
rect 170 10 172 12
rect 174 10 176 12
rect 170 8 176 10
rect 210 12 216 14
rect 210 10 212 12
rect 214 10 216 12
rect 210 8 216 10
rect 309 12 315 14
rect 309 10 311 12
rect 313 10 315 12
rect 309 8 315 10
rect 523 12 529 14
rect 523 10 525 12
rect 527 10 529 12
rect 523 8 529 10
rect 617 12 623 14
rect 617 10 619 12
rect 621 10 623 12
rect 617 8 623 10
<< ntie >>
rect 7 516 13 518
rect 7 514 9 516
rect 11 514 13 516
rect 56 516 62 518
rect 7 512 13 514
rect 56 514 58 516
rect 60 514 62 516
rect 129 516 135 518
rect 56 512 62 514
rect 129 514 131 516
rect 133 514 135 516
rect 170 516 176 518
rect 129 512 135 514
rect 170 514 172 516
rect 174 514 176 516
rect 243 516 249 518
rect 170 512 176 514
rect 243 514 245 516
rect 247 514 249 516
rect 309 516 315 518
rect 243 512 249 514
rect 309 514 311 516
rect 313 514 315 516
rect 523 516 529 518
rect 309 512 315 514
rect 523 514 525 516
rect 527 514 529 516
rect 584 516 590 518
rect 523 512 529 514
rect 584 514 586 516
rect 588 514 590 516
rect 584 512 590 514
rect 7 504 13 506
rect 7 502 9 504
rect 11 502 13 504
rect 56 504 62 506
rect 7 500 13 502
rect 56 502 58 504
rect 60 502 62 504
rect 129 504 135 506
rect 56 500 62 502
rect 129 502 131 504
rect 133 502 135 504
rect 170 504 176 506
rect 129 500 135 502
rect 170 502 172 504
rect 174 502 176 504
rect 243 504 249 506
rect 170 500 176 502
rect 243 502 245 504
rect 247 502 249 504
rect 309 504 315 506
rect 243 500 249 502
rect 309 502 311 504
rect 313 502 315 504
rect 523 504 529 506
rect 309 500 315 502
rect 523 502 525 504
rect 527 502 529 504
rect 584 504 590 506
rect 523 500 529 502
rect 584 502 586 504
rect 588 502 590 504
rect 584 500 590 502
rect 7 372 13 374
rect 7 370 9 372
rect 11 370 13 372
rect 56 372 62 374
rect 7 368 13 370
rect 56 370 58 372
rect 60 370 62 372
rect 129 372 135 374
rect 56 368 62 370
rect 129 370 131 372
rect 133 370 135 372
rect 170 372 176 374
rect 129 368 135 370
rect 170 370 172 372
rect 174 370 176 372
rect 243 372 249 374
rect 170 368 176 370
rect 243 370 245 372
rect 247 370 249 372
rect 309 372 315 374
rect 243 368 249 370
rect 309 370 311 372
rect 313 370 315 372
rect 523 372 529 374
rect 309 368 315 370
rect 523 370 525 372
rect 527 370 529 372
rect 584 372 590 374
rect 523 368 529 370
rect 584 370 586 372
rect 588 370 590 372
rect 584 368 590 370
rect 7 360 13 362
rect 7 358 9 360
rect 11 358 13 360
rect 56 360 62 362
rect 7 356 13 358
rect 56 358 58 360
rect 60 358 62 360
rect 129 360 135 362
rect 56 356 62 358
rect 129 358 131 360
rect 133 358 135 360
rect 170 360 176 362
rect 129 356 135 358
rect 170 358 172 360
rect 174 358 176 360
rect 243 360 249 362
rect 170 356 176 358
rect 243 358 245 360
rect 247 358 249 360
rect 309 360 315 362
rect 243 356 249 358
rect 309 358 311 360
rect 313 358 315 360
rect 523 360 529 362
rect 309 356 315 358
rect 523 358 525 360
rect 527 358 529 360
rect 584 360 590 362
rect 523 356 529 358
rect 584 358 586 360
rect 588 358 590 360
rect 584 356 590 358
rect 7 228 13 230
rect 7 226 9 228
rect 11 226 13 228
rect 56 228 62 230
rect 7 224 13 226
rect 56 226 58 228
rect 60 226 62 228
rect 129 228 135 230
rect 56 224 62 226
rect 129 226 131 228
rect 133 226 135 228
rect 170 228 176 230
rect 129 224 135 226
rect 170 226 172 228
rect 174 226 176 228
rect 243 228 249 230
rect 170 224 176 226
rect 243 226 245 228
rect 247 226 249 228
rect 309 228 315 230
rect 243 224 249 226
rect 309 226 311 228
rect 313 226 315 228
rect 523 228 529 230
rect 309 224 315 226
rect 523 226 525 228
rect 527 226 529 228
rect 584 228 590 230
rect 523 224 529 226
rect 584 226 586 228
rect 588 226 590 228
rect 584 224 590 226
rect 7 216 13 218
rect 7 214 9 216
rect 11 214 13 216
rect 56 216 62 218
rect 7 212 13 214
rect 56 214 58 216
rect 60 214 62 216
rect 129 216 135 218
rect 56 212 62 214
rect 129 214 131 216
rect 133 214 135 216
rect 170 216 176 218
rect 129 212 135 214
rect 170 214 172 216
rect 174 214 176 216
rect 243 216 249 218
rect 170 212 176 214
rect 243 214 245 216
rect 247 214 249 216
rect 309 216 315 218
rect 243 212 249 214
rect 309 214 311 216
rect 313 214 315 216
rect 523 216 529 218
rect 309 212 315 214
rect 523 214 525 216
rect 527 214 529 216
rect 584 216 590 218
rect 523 212 529 214
rect 584 214 586 216
rect 588 214 590 216
rect 584 212 590 214
rect 7 84 13 86
rect 7 82 9 84
rect 11 82 13 84
rect 56 84 62 86
rect 7 80 13 82
rect 56 82 58 84
rect 60 82 62 84
rect 129 84 135 86
rect 56 80 62 82
rect 129 82 131 84
rect 133 82 135 84
rect 170 84 176 86
rect 129 80 135 82
rect 170 82 172 84
rect 174 82 176 84
rect 243 84 249 86
rect 170 80 176 82
rect 243 82 245 84
rect 247 82 249 84
rect 309 84 315 86
rect 243 80 249 82
rect 309 82 311 84
rect 313 82 315 84
rect 523 84 529 86
rect 309 80 315 82
rect 523 82 525 84
rect 527 82 529 84
rect 584 84 590 86
rect 523 80 529 82
rect 584 82 586 84
rect 588 82 590 84
rect 584 80 590 82
rect 7 72 13 74
rect 7 70 9 72
rect 11 70 13 72
rect 56 72 62 74
rect 7 68 13 70
rect 56 70 58 72
rect 60 70 62 72
rect 129 72 135 74
rect 56 68 62 70
rect 129 70 131 72
rect 133 70 135 72
rect 170 72 176 74
rect 129 68 135 70
rect 170 70 172 72
rect 174 70 176 72
rect 243 72 249 74
rect 170 68 176 70
rect 243 70 245 72
rect 247 70 249 72
rect 309 72 315 74
rect 243 68 249 70
rect 309 70 311 72
rect 313 70 315 72
rect 523 72 529 74
rect 309 68 315 70
rect 523 70 525 72
rect 527 70 529 72
rect 584 72 590 74
rect 523 68 529 70
rect 584 70 586 72
rect 588 70 590 72
rect 584 68 590 70
<< nmos >>
rect 13 555 15 564
rect 23 555 25 561
rect 33 555 35 561
rect 62 557 64 566
rect 75 557 77 568
rect 82 557 84 568
rect 102 555 104 564
rect 118 560 120 569
rect 128 560 130 569
rect 138 560 140 572
rect 145 560 147 572
rect 176 557 178 566
rect 189 557 191 568
rect 196 557 198 568
rect 216 555 218 564
rect 232 560 234 569
rect 242 560 244 569
rect 252 560 254 572
rect 259 560 261 572
rect 287 557 289 568
rect 294 557 296 568
rect 307 557 309 566
rect 329 561 331 567
rect 339 561 341 569
rect 346 561 348 569
rect 356 561 358 569
rect 363 561 365 569
rect 373 560 375 569
rect 396 560 398 569
rect 406 561 408 569
rect 413 561 415 569
rect 423 561 425 569
rect 430 561 432 569
rect 440 561 442 567
rect 463 560 465 569
rect 473 561 475 569
rect 480 561 482 569
rect 490 561 492 569
rect 497 561 499 569
rect 507 561 509 567
rect 529 555 531 564
rect 539 555 541 561
rect 549 555 551 561
rect 572 560 574 572
rect 579 560 581 572
rect 589 560 591 569
rect 599 560 601 569
rect 615 555 617 564
rect 13 454 15 463
rect 23 457 25 463
rect 33 457 35 463
rect 62 452 64 461
rect 75 450 77 461
rect 82 450 84 461
rect 102 454 104 463
rect 118 449 120 458
rect 128 449 130 458
rect 138 446 140 458
rect 145 446 147 458
rect 176 452 178 461
rect 189 450 191 461
rect 196 450 198 461
rect 216 454 218 463
rect 232 449 234 458
rect 242 449 244 458
rect 252 446 254 458
rect 259 446 261 458
rect 287 450 289 461
rect 294 450 296 461
rect 307 452 309 461
rect 329 451 331 457
rect 339 449 341 457
rect 346 449 348 457
rect 356 449 358 457
rect 363 449 365 457
rect 373 449 375 458
rect 396 449 398 458
rect 406 449 408 457
rect 413 449 415 457
rect 423 449 425 457
rect 430 449 432 457
rect 440 451 442 457
rect 463 449 465 458
rect 473 449 475 457
rect 480 449 482 457
rect 490 449 492 457
rect 497 449 499 457
rect 507 451 509 457
rect 529 454 531 463
rect 539 457 541 463
rect 549 457 551 463
rect 572 446 574 458
rect 579 446 581 458
rect 589 449 591 458
rect 599 449 601 458
rect 615 454 617 463
rect 13 411 15 420
rect 23 411 25 417
rect 33 411 35 417
rect 62 413 64 422
rect 75 413 77 424
rect 82 413 84 424
rect 102 411 104 420
rect 118 416 120 425
rect 128 416 130 425
rect 138 416 140 428
rect 145 416 147 428
rect 176 413 178 422
rect 189 413 191 424
rect 196 413 198 424
rect 216 411 218 420
rect 232 416 234 425
rect 242 416 244 425
rect 252 416 254 428
rect 259 416 261 428
rect 287 413 289 424
rect 294 413 296 424
rect 307 413 309 422
rect 329 417 331 423
rect 339 417 341 425
rect 346 417 348 425
rect 356 417 358 425
rect 363 417 365 425
rect 373 416 375 425
rect 396 416 398 425
rect 406 417 408 425
rect 413 417 415 425
rect 423 417 425 425
rect 430 417 432 425
rect 440 417 442 423
rect 463 416 465 425
rect 473 417 475 425
rect 480 417 482 425
rect 490 417 492 425
rect 497 417 499 425
rect 507 417 509 423
rect 529 411 531 420
rect 539 411 541 417
rect 549 411 551 417
rect 572 416 574 428
rect 579 416 581 428
rect 589 416 591 425
rect 599 416 601 425
rect 615 411 617 420
rect 13 310 15 319
rect 23 313 25 319
rect 33 313 35 319
rect 62 308 64 317
rect 75 306 77 317
rect 82 306 84 317
rect 102 310 104 319
rect 118 305 120 314
rect 128 305 130 314
rect 138 302 140 314
rect 145 302 147 314
rect 176 308 178 317
rect 189 306 191 317
rect 196 306 198 317
rect 216 310 218 319
rect 232 305 234 314
rect 242 305 244 314
rect 252 302 254 314
rect 259 302 261 314
rect 287 306 289 317
rect 294 306 296 317
rect 307 308 309 317
rect 329 307 331 313
rect 339 305 341 313
rect 346 305 348 313
rect 356 305 358 313
rect 363 305 365 313
rect 373 305 375 314
rect 396 305 398 314
rect 406 305 408 313
rect 413 305 415 313
rect 423 305 425 313
rect 430 305 432 313
rect 440 307 442 313
rect 463 305 465 314
rect 473 305 475 313
rect 480 305 482 313
rect 490 305 492 313
rect 497 305 499 313
rect 507 307 509 313
rect 529 310 531 319
rect 539 313 541 319
rect 549 313 551 319
rect 572 302 574 314
rect 579 302 581 314
rect 589 305 591 314
rect 599 305 601 314
rect 615 310 617 319
rect 13 267 15 276
rect 23 267 25 273
rect 33 267 35 273
rect 62 269 64 278
rect 75 269 77 280
rect 82 269 84 280
rect 102 267 104 276
rect 118 272 120 281
rect 128 272 130 281
rect 138 272 140 284
rect 145 272 147 284
rect 176 269 178 278
rect 189 269 191 280
rect 196 269 198 280
rect 216 267 218 276
rect 232 272 234 281
rect 242 272 244 281
rect 252 272 254 284
rect 259 272 261 284
rect 287 269 289 280
rect 294 269 296 280
rect 307 269 309 278
rect 329 273 331 279
rect 339 273 341 281
rect 346 273 348 281
rect 356 273 358 281
rect 363 273 365 281
rect 373 272 375 281
rect 396 272 398 281
rect 406 273 408 281
rect 413 273 415 281
rect 423 273 425 281
rect 430 273 432 281
rect 440 273 442 279
rect 463 272 465 281
rect 473 273 475 281
rect 480 273 482 281
rect 490 273 492 281
rect 497 273 499 281
rect 507 273 509 279
rect 529 267 531 276
rect 539 267 541 273
rect 549 267 551 273
rect 572 272 574 284
rect 579 272 581 284
rect 589 272 591 281
rect 599 272 601 281
rect 615 267 617 276
rect 13 166 15 175
rect 23 169 25 175
rect 33 169 35 175
rect 62 164 64 173
rect 75 162 77 173
rect 82 162 84 173
rect 102 166 104 175
rect 118 161 120 170
rect 128 161 130 170
rect 138 158 140 170
rect 145 158 147 170
rect 176 164 178 173
rect 189 162 191 173
rect 196 162 198 173
rect 216 166 218 175
rect 232 161 234 170
rect 242 161 244 170
rect 252 158 254 170
rect 259 158 261 170
rect 287 162 289 173
rect 294 162 296 173
rect 307 164 309 173
rect 329 163 331 169
rect 339 161 341 169
rect 346 161 348 169
rect 356 161 358 169
rect 363 161 365 169
rect 373 161 375 170
rect 396 161 398 170
rect 406 161 408 169
rect 413 161 415 169
rect 423 161 425 169
rect 430 161 432 169
rect 440 163 442 169
rect 463 161 465 170
rect 473 161 475 169
rect 480 161 482 169
rect 490 161 492 169
rect 497 161 499 169
rect 507 163 509 169
rect 529 166 531 175
rect 539 169 541 175
rect 549 169 551 175
rect 572 158 574 170
rect 579 158 581 170
rect 589 161 591 170
rect 599 161 601 170
rect 615 166 617 175
rect 13 123 15 132
rect 23 123 25 129
rect 33 123 35 129
rect 62 125 64 134
rect 75 125 77 136
rect 82 125 84 136
rect 102 123 104 132
rect 118 128 120 137
rect 128 128 130 137
rect 138 128 140 140
rect 145 128 147 140
rect 176 125 178 134
rect 189 125 191 136
rect 196 125 198 136
rect 216 123 218 132
rect 232 128 234 137
rect 242 128 244 137
rect 252 128 254 140
rect 259 128 261 140
rect 287 125 289 136
rect 294 125 296 136
rect 307 125 309 134
rect 329 129 331 135
rect 339 129 341 137
rect 346 129 348 137
rect 356 129 358 137
rect 363 129 365 137
rect 373 128 375 137
rect 396 128 398 137
rect 406 129 408 137
rect 413 129 415 137
rect 423 129 425 137
rect 430 129 432 137
rect 440 129 442 135
rect 463 128 465 137
rect 473 129 475 137
rect 480 129 482 137
rect 490 129 492 137
rect 497 129 499 137
rect 507 129 509 135
rect 529 123 531 132
rect 539 123 541 129
rect 549 123 551 129
rect 572 128 574 140
rect 579 128 581 140
rect 589 128 591 137
rect 599 128 601 137
rect 615 123 617 132
rect 13 22 15 31
rect 23 25 25 31
rect 33 25 35 31
rect 62 20 64 29
rect 75 18 77 29
rect 82 18 84 29
rect 102 22 104 31
rect 118 17 120 26
rect 128 17 130 26
rect 138 14 140 26
rect 145 14 147 26
rect 176 20 178 29
rect 189 18 191 29
rect 196 18 198 29
rect 216 22 218 31
rect 232 17 234 26
rect 242 17 244 26
rect 252 14 254 26
rect 259 14 261 26
rect 287 18 289 29
rect 294 18 296 29
rect 307 20 309 29
rect 329 19 331 25
rect 339 17 341 25
rect 346 17 348 25
rect 356 17 358 25
rect 363 17 365 25
rect 373 17 375 26
rect 396 17 398 26
rect 406 17 408 25
rect 413 17 415 25
rect 423 17 425 25
rect 430 17 432 25
rect 440 19 442 25
rect 463 17 465 26
rect 473 17 475 25
rect 480 17 482 25
rect 490 17 492 25
rect 497 17 499 25
rect 507 19 509 25
rect 529 22 531 31
rect 539 25 541 31
rect 549 25 551 31
rect 572 14 574 26
rect 579 14 581 26
rect 589 17 591 26
rect 599 17 601 26
rect 615 22 617 31
<< pmos >>
rect 13 525 15 543
rect 26 515 28 536
rect 33 515 35 536
rect 62 524 64 542
rect 72 522 74 535
rect 82 522 84 535
rect 110 515 112 542
rect 126 524 128 542
rect 136 524 138 542
rect 146 515 148 542
rect 176 524 178 542
rect 186 522 188 535
rect 196 522 198 535
rect 224 515 226 542
rect 240 524 242 542
rect 250 524 252 542
rect 260 515 262 542
rect 287 522 289 535
rect 297 522 299 535
rect 307 524 309 542
rect 329 535 331 543
rect 339 515 341 531
rect 346 515 348 531
rect 356 515 358 531
rect 363 515 365 531
rect 373 515 375 533
rect 396 515 398 533
rect 440 535 442 543
rect 406 515 408 531
rect 413 515 415 531
rect 423 515 425 531
rect 430 515 432 531
rect 463 515 465 533
rect 507 535 509 543
rect 473 515 475 531
rect 480 515 482 531
rect 490 515 492 531
rect 497 515 499 531
rect 529 525 531 543
rect 542 515 544 536
rect 549 515 551 536
rect 571 515 573 542
rect 581 524 583 542
rect 591 524 593 542
rect 607 515 609 542
rect 13 475 15 493
rect 26 482 28 503
rect 33 482 35 503
rect 62 476 64 494
rect 72 483 74 496
rect 82 483 84 496
rect 110 476 112 503
rect 126 476 128 494
rect 136 476 138 494
rect 146 476 148 503
rect 176 476 178 494
rect 186 483 188 496
rect 196 483 198 496
rect 224 476 226 503
rect 240 476 242 494
rect 250 476 252 494
rect 260 476 262 503
rect 287 483 289 496
rect 297 483 299 496
rect 307 476 309 494
rect 339 487 341 503
rect 346 487 348 503
rect 356 487 358 503
rect 363 487 365 503
rect 329 475 331 483
rect 373 485 375 503
rect 396 485 398 503
rect 406 487 408 503
rect 413 487 415 503
rect 423 487 425 503
rect 430 487 432 503
rect 463 485 465 503
rect 473 487 475 503
rect 480 487 482 503
rect 490 487 492 503
rect 497 487 499 503
rect 440 475 442 483
rect 507 475 509 483
rect 529 475 531 493
rect 542 482 544 503
rect 549 482 551 503
rect 571 476 573 503
rect 581 476 583 494
rect 591 476 593 494
rect 607 476 609 503
rect 13 381 15 399
rect 26 371 28 392
rect 33 371 35 392
rect 62 380 64 398
rect 72 378 74 391
rect 82 378 84 391
rect 110 371 112 398
rect 126 380 128 398
rect 136 380 138 398
rect 146 371 148 398
rect 176 380 178 398
rect 186 378 188 391
rect 196 378 198 391
rect 224 371 226 398
rect 240 380 242 398
rect 250 380 252 398
rect 260 371 262 398
rect 287 378 289 391
rect 297 378 299 391
rect 307 380 309 398
rect 329 391 331 399
rect 339 371 341 387
rect 346 371 348 387
rect 356 371 358 387
rect 363 371 365 387
rect 373 371 375 389
rect 396 371 398 389
rect 440 391 442 399
rect 406 371 408 387
rect 413 371 415 387
rect 423 371 425 387
rect 430 371 432 387
rect 463 371 465 389
rect 507 391 509 399
rect 473 371 475 387
rect 480 371 482 387
rect 490 371 492 387
rect 497 371 499 387
rect 529 381 531 399
rect 542 371 544 392
rect 549 371 551 392
rect 571 371 573 398
rect 581 380 583 398
rect 591 380 593 398
rect 607 371 609 398
rect 13 331 15 349
rect 26 338 28 359
rect 33 338 35 359
rect 62 332 64 350
rect 72 339 74 352
rect 82 339 84 352
rect 110 332 112 359
rect 126 332 128 350
rect 136 332 138 350
rect 146 332 148 359
rect 176 332 178 350
rect 186 339 188 352
rect 196 339 198 352
rect 224 332 226 359
rect 240 332 242 350
rect 250 332 252 350
rect 260 332 262 359
rect 287 339 289 352
rect 297 339 299 352
rect 307 332 309 350
rect 339 343 341 359
rect 346 343 348 359
rect 356 343 358 359
rect 363 343 365 359
rect 329 331 331 339
rect 373 341 375 359
rect 396 341 398 359
rect 406 343 408 359
rect 413 343 415 359
rect 423 343 425 359
rect 430 343 432 359
rect 463 341 465 359
rect 473 343 475 359
rect 480 343 482 359
rect 490 343 492 359
rect 497 343 499 359
rect 440 331 442 339
rect 507 331 509 339
rect 529 331 531 349
rect 542 338 544 359
rect 549 338 551 359
rect 571 332 573 359
rect 581 332 583 350
rect 591 332 593 350
rect 607 332 609 359
rect 13 237 15 255
rect 26 227 28 248
rect 33 227 35 248
rect 62 236 64 254
rect 72 234 74 247
rect 82 234 84 247
rect 110 227 112 254
rect 126 236 128 254
rect 136 236 138 254
rect 146 227 148 254
rect 176 236 178 254
rect 186 234 188 247
rect 196 234 198 247
rect 224 227 226 254
rect 240 236 242 254
rect 250 236 252 254
rect 260 227 262 254
rect 287 234 289 247
rect 297 234 299 247
rect 307 236 309 254
rect 329 247 331 255
rect 339 227 341 243
rect 346 227 348 243
rect 356 227 358 243
rect 363 227 365 243
rect 373 227 375 245
rect 396 227 398 245
rect 440 247 442 255
rect 406 227 408 243
rect 413 227 415 243
rect 423 227 425 243
rect 430 227 432 243
rect 463 227 465 245
rect 507 247 509 255
rect 473 227 475 243
rect 480 227 482 243
rect 490 227 492 243
rect 497 227 499 243
rect 529 237 531 255
rect 542 227 544 248
rect 549 227 551 248
rect 571 227 573 254
rect 581 236 583 254
rect 591 236 593 254
rect 607 227 609 254
rect 13 187 15 205
rect 26 194 28 215
rect 33 194 35 215
rect 62 188 64 206
rect 72 195 74 208
rect 82 195 84 208
rect 110 188 112 215
rect 126 188 128 206
rect 136 188 138 206
rect 146 188 148 215
rect 176 188 178 206
rect 186 195 188 208
rect 196 195 198 208
rect 224 188 226 215
rect 240 188 242 206
rect 250 188 252 206
rect 260 188 262 215
rect 287 195 289 208
rect 297 195 299 208
rect 307 188 309 206
rect 339 199 341 215
rect 346 199 348 215
rect 356 199 358 215
rect 363 199 365 215
rect 329 187 331 195
rect 373 197 375 215
rect 396 197 398 215
rect 406 199 408 215
rect 413 199 415 215
rect 423 199 425 215
rect 430 199 432 215
rect 463 197 465 215
rect 473 199 475 215
rect 480 199 482 215
rect 490 199 492 215
rect 497 199 499 215
rect 440 187 442 195
rect 507 187 509 195
rect 529 187 531 205
rect 542 194 544 215
rect 549 194 551 215
rect 571 188 573 215
rect 581 188 583 206
rect 591 188 593 206
rect 607 188 609 215
rect 13 93 15 111
rect 26 83 28 104
rect 33 83 35 104
rect 62 92 64 110
rect 72 90 74 103
rect 82 90 84 103
rect 110 83 112 110
rect 126 92 128 110
rect 136 92 138 110
rect 146 83 148 110
rect 176 92 178 110
rect 186 90 188 103
rect 196 90 198 103
rect 224 83 226 110
rect 240 92 242 110
rect 250 92 252 110
rect 260 83 262 110
rect 287 90 289 103
rect 297 90 299 103
rect 307 92 309 110
rect 329 103 331 111
rect 339 83 341 99
rect 346 83 348 99
rect 356 83 358 99
rect 363 83 365 99
rect 373 83 375 101
rect 396 83 398 101
rect 440 103 442 111
rect 406 83 408 99
rect 413 83 415 99
rect 423 83 425 99
rect 430 83 432 99
rect 463 83 465 101
rect 507 103 509 111
rect 473 83 475 99
rect 480 83 482 99
rect 490 83 492 99
rect 497 83 499 99
rect 529 93 531 111
rect 542 83 544 104
rect 549 83 551 104
rect 571 83 573 110
rect 581 92 583 110
rect 591 92 593 110
rect 607 83 609 110
rect 13 43 15 61
rect 26 50 28 71
rect 33 50 35 71
rect 62 44 64 62
rect 72 51 74 64
rect 82 51 84 64
rect 110 44 112 71
rect 126 44 128 62
rect 136 44 138 62
rect 146 44 148 71
rect 176 44 178 62
rect 186 51 188 64
rect 196 51 198 64
rect 224 44 226 71
rect 240 44 242 62
rect 250 44 252 62
rect 260 44 262 71
rect 287 51 289 64
rect 297 51 299 64
rect 307 44 309 62
rect 339 55 341 71
rect 346 55 348 71
rect 356 55 358 71
rect 363 55 365 71
rect 329 43 331 51
rect 373 53 375 71
rect 396 53 398 71
rect 406 55 408 71
rect 413 55 415 71
rect 423 55 425 71
rect 430 55 432 71
rect 463 53 465 71
rect 473 55 475 71
rect 480 55 482 71
rect 490 55 492 71
rect 497 55 499 71
rect 440 43 442 51
rect 507 43 509 51
rect 529 43 531 61
rect 542 50 544 71
rect 549 50 551 71
rect 571 44 573 71
rect 581 44 583 62
rect 591 44 593 62
rect 607 44 609 71
<< polyct0 >>
rect 15 548 17 550
rect 64 548 66 550
rect 134 548 136 550
rect 144 547 146 549
rect 178 548 180 550
rect 248 548 250 550
rect 258 547 260 549
rect 305 548 307 550
rect 354 554 356 556
rect 372 553 374 555
rect 397 553 399 555
rect 347 538 349 540
rect 415 554 417 556
rect 422 538 424 540
rect 464 553 466 555
rect 482 554 484 556
rect 489 538 491 540
rect 531 548 533 550
rect 573 547 575 549
rect 583 548 585 550
rect 15 468 17 470
rect 64 468 66 470
rect 134 468 136 470
rect 144 469 146 471
rect 178 468 180 470
rect 248 468 250 470
rect 258 469 260 471
rect 305 468 307 470
rect 347 478 349 480
rect 354 462 356 464
rect 422 478 424 480
rect 372 463 374 465
rect 397 463 399 465
rect 415 462 417 464
rect 489 478 491 480
rect 464 463 466 465
rect 482 462 484 464
rect 531 468 533 470
rect 573 469 575 471
rect 583 468 585 470
rect 15 404 17 406
rect 64 404 66 406
rect 134 404 136 406
rect 144 403 146 405
rect 178 404 180 406
rect 248 404 250 406
rect 258 403 260 405
rect 305 404 307 406
rect 354 410 356 412
rect 372 409 374 411
rect 397 409 399 411
rect 347 394 349 396
rect 415 410 417 412
rect 422 394 424 396
rect 464 409 466 411
rect 482 410 484 412
rect 489 394 491 396
rect 531 404 533 406
rect 573 403 575 405
rect 583 404 585 406
rect 15 324 17 326
rect 64 324 66 326
rect 134 324 136 326
rect 144 325 146 327
rect 178 324 180 326
rect 248 324 250 326
rect 258 325 260 327
rect 305 324 307 326
rect 347 334 349 336
rect 354 318 356 320
rect 422 334 424 336
rect 372 319 374 321
rect 397 319 399 321
rect 415 318 417 320
rect 489 334 491 336
rect 464 319 466 321
rect 482 318 484 320
rect 531 324 533 326
rect 573 325 575 327
rect 583 324 585 326
rect 15 260 17 262
rect 64 260 66 262
rect 134 260 136 262
rect 144 259 146 261
rect 178 260 180 262
rect 248 260 250 262
rect 258 259 260 261
rect 305 260 307 262
rect 354 266 356 268
rect 372 265 374 267
rect 397 265 399 267
rect 347 250 349 252
rect 415 266 417 268
rect 422 250 424 252
rect 464 265 466 267
rect 482 266 484 268
rect 489 250 491 252
rect 531 260 533 262
rect 573 259 575 261
rect 583 260 585 262
rect 15 180 17 182
rect 64 180 66 182
rect 134 180 136 182
rect 144 181 146 183
rect 178 180 180 182
rect 248 180 250 182
rect 258 181 260 183
rect 305 180 307 182
rect 347 190 349 192
rect 354 174 356 176
rect 422 190 424 192
rect 372 175 374 177
rect 397 175 399 177
rect 415 174 417 176
rect 489 190 491 192
rect 464 175 466 177
rect 482 174 484 176
rect 531 180 533 182
rect 573 181 575 183
rect 583 180 585 182
rect 15 116 17 118
rect 64 116 66 118
rect 134 116 136 118
rect 144 115 146 117
rect 178 116 180 118
rect 248 116 250 118
rect 258 115 260 117
rect 305 116 307 118
rect 354 122 356 124
rect 372 121 374 123
rect 397 121 399 123
rect 347 106 349 108
rect 415 122 417 124
rect 422 106 424 108
rect 464 121 466 123
rect 482 122 484 124
rect 489 106 491 108
rect 531 116 533 118
rect 573 115 575 117
rect 583 116 585 118
rect 15 36 17 38
rect 64 36 66 38
rect 134 36 136 38
rect 144 37 146 39
rect 178 36 180 38
rect 248 36 250 38
rect 258 37 260 39
rect 305 36 307 38
rect 347 46 349 48
rect 354 30 356 32
rect 422 46 424 48
rect 372 31 374 33
rect 397 31 399 33
rect 415 30 417 32
rect 489 46 491 48
rect 464 31 466 33
rect 482 30 484 32
rect 531 36 533 38
rect 573 37 575 39
rect 583 36 585 38
<< polyct1 >>
rect 25 548 27 550
rect 74 548 76 550
rect 35 541 37 543
rect 113 553 115 555
rect 84 540 86 542
rect 188 548 190 550
rect 97 540 99 542
rect 227 553 229 555
rect 198 540 200 542
rect 295 548 297 550
rect 211 540 213 542
rect 285 540 287 542
rect 337 548 339 550
rect 364 543 366 545
rect 405 543 407 545
rect 432 548 434 550
rect 324 528 326 530
rect 472 543 474 545
rect 499 548 501 550
rect 445 528 447 530
rect 541 548 543 550
rect 512 528 514 530
rect 604 553 606 555
rect 551 541 553 543
rect 620 540 622 542
rect 35 475 37 477
rect 25 468 27 470
rect 84 476 86 478
rect 97 476 99 478
rect 74 468 76 470
rect 198 476 200 478
rect 211 476 213 478
rect 285 476 287 478
rect 113 463 115 465
rect 188 468 190 470
rect 227 463 229 465
rect 324 488 326 490
rect 295 468 297 470
rect 445 488 447 490
rect 337 468 339 470
rect 364 473 366 475
rect 405 473 407 475
rect 512 488 514 490
rect 432 468 434 470
rect 472 473 474 475
rect 499 468 501 470
rect 551 475 553 477
rect 620 476 622 478
rect 541 468 543 470
rect 604 463 606 465
rect 25 404 27 406
rect 74 404 76 406
rect 35 397 37 399
rect 113 409 115 411
rect 84 396 86 398
rect 188 404 190 406
rect 97 396 99 398
rect 227 409 229 411
rect 198 396 200 398
rect 295 404 297 406
rect 211 396 213 398
rect 285 396 287 398
rect 337 404 339 406
rect 364 399 366 401
rect 405 399 407 401
rect 432 404 434 406
rect 324 384 326 386
rect 472 399 474 401
rect 499 404 501 406
rect 445 384 447 386
rect 541 404 543 406
rect 512 384 514 386
rect 604 409 606 411
rect 551 397 553 399
rect 620 396 622 398
rect 35 331 37 333
rect 25 324 27 326
rect 84 332 86 334
rect 97 332 99 334
rect 74 324 76 326
rect 198 332 200 334
rect 211 332 213 334
rect 285 332 287 334
rect 113 319 115 321
rect 188 324 190 326
rect 227 319 229 321
rect 324 344 326 346
rect 295 324 297 326
rect 445 344 447 346
rect 337 324 339 326
rect 364 329 366 331
rect 405 329 407 331
rect 512 344 514 346
rect 432 324 434 326
rect 472 329 474 331
rect 499 324 501 326
rect 551 331 553 333
rect 620 332 622 334
rect 541 324 543 326
rect 604 319 606 321
rect 25 260 27 262
rect 74 260 76 262
rect 35 253 37 255
rect 113 265 115 267
rect 84 252 86 254
rect 188 260 190 262
rect 97 252 99 254
rect 227 265 229 267
rect 198 252 200 254
rect 295 260 297 262
rect 211 252 213 254
rect 285 252 287 254
rect 337 260 339 262
rect 364 255 366 257
rect 405 255 407 257
rect 432 260 434 262
rect 324 240 326 242
rect 472 255 474 257
rect 499 260 501 262
rect 445 240 447 242
rect 541 260 543 262
rect 512 240 514 242
rect 604 265 606 267
rect 551 253 553 255
rect 620 252 622 254
rect 35 187 37 189
rect 25 180 27 182
rect 84 188 86 190
rect 97 188 99 190
rect 74 180 76 182
rect 198 188 200 190
rect 211 188 213 190
rect 285 188 287 190
rect 113 175 115 177
rect 188 180 190 182
rect 227 175 229 177
rect 324 200 326 202
rect 295 180 297 182
rect 445 200 447 202
rect 337 180 339 182
rect 364 185 366 187
rect 405 185 407 187
rect 512 200 514 202
rect 432 180 434 182
rect 472 185 474 187
rect 499 180 501 182
rect 551 187 553 189
rect 620 188 622 190
rect 541 180 543 182
rect 604 175 606 177
rect 25 116 27 118
rect 74 116 76 118
rect 35 109 37 111
rect 113 121 115 123
rect 84 108 86 110
rect 188 116 190 118
rect 97 108 99 110
rect 227 121 229 123
rect 198 108 200 110
rect 295 116 297 118
rect 211 108 213 110
rect 285 108 287 110
rect 337 116 339 118
rect 364 111 366 113
rect 405 111 407 113
rect 432 116 434 118
rect 324 96 326 98
rect 472 111 474 113
rect 499 116 501 118
rect 445 96 447 98
rect 541 116 543 118
rect 512 96 514 98
rect 604 121 606 123
rect 551 109 553 111
rect 620 108 622 110
rect 35 43 37 45
rect 25 36 27 38
rect 84 44 86 46
rect 97 44 99 46
rect 74 36 76 38
rect 198 44 200 46
rect 211 44 213 46
rect 285 44 287 46
rect 113 31 115 33
rect 188 36 190 38
rect 227 31 229 33
rect 324 56 326 58
rect 295 36 297 38
rect 445 56 447 58
rect 337 36 339 38
rect 364 41 366 43
rect 405 41 407 43
rect 512 56 514 58
rect 432 36 434 38
rect 472 41 474 43
rect 499 36 501 38
rect 551 43 553 45
rect 620 44 622 46
rect 541 36 543 38
rect 604 31 606 33
<< ndifct0 >>
rect 19 570 21 572
rect 38 570 40 572
rect 28 557 30 559
rect 87 564 89 566
rect 111 565 113 567
rect 97 557 99 559
rect 123 562 125 564
rect 201 564 203 566
rect 225 565 227 567
rect 211 557 213 559
rect 237 562 239 564
rect 282 564 284 566
rect 324 563 326 565
rect 334 563 336 565
rect 351 565 353 567
rect 368 565 370 567
rect 401 565 403 567
rect 418 565 420 567
rect 435 563 437 565
rect 445 563 447 565
rect 468 565 470 567
rect 485 565 487 567
rect 535 570 537 572
rect 502 563 504 565
rect 512 563 514 565
rect 554 570 556 572
rect 544 557 546 559
rect 594 562 596 564
rect 606 565 608 567
rect 620 557 622 559
rect 28 459 30 461
rect 19 446 21 448
rect 97 459 99 461
rect 87 452 89 454
rect 111 451 113 453
rect 38 446 40 448
rect 123 454 125 456
rect 211 459 213 461
rect 201 452 203 454
rect 225 451 227 453
rect 237 454 239 456
rect 282 452 284 454
rect 324 453 326 455
rect 334 453 336 455
rect 351 451 353 453
rect 368 451 370 453
rect 401 451 403 453
rect 418 451 420 453
rect 435 453 437 455
rect 445 453 447 455
rect 468 451 470 453
rect 485 451 487 453
rect 502 453 504 455
rect 512 453 514 455
rect 544 459 546 461
rect 535 446 537 448
rect 554 446 556 448
rect 594 454 596 456
rect 620 459 622 461
rect 606 451 608 453
rect 19 426 21 428
rect 38 426 40 428
rect 28 413 30 415
rect 87 420 89 422
rect 111 421 113 423
rect 97 413 99 415
rect 123 418 125 420
rect 201 420 203 422
rect 225 421 227 423
rect 211 413 213 415
rect 237 418 239 420
rect 282 420 284 422
rect 324 419 326 421
rect 334 419 336 421
rect 351 421 353 423
rect 368 421 370 423
rect 401 421 403 423
rect 418 421 420 423
rect 435 419 437 421
rect 445 419 447 421
rect 468 421 470 423
rect 485 421 487 423
rect 535 426 537 428
rect 502 419 504 421
rect 512 419 514 421
rect 554 426 556 428
rect 544 413 546 415
rect 594 418 596 420
rect 606 421 608 423
rect 620 413 622 415
rect 28 315 30 317
rect 19 302 21 304
rect 97 315 99 317
rect 87 308 89 310
rect 111 307 113 309
rect 38 302 40 304
rect 123 310 125 312
rect 211 315 213 317
rect 201 308 203 310
rect 225 307 227 309
rect 237 310 239 312
rect 282 308 284 310
rect 324 309 326 311
rect 334 309 336 311
rect 351 307 353 309
rect 368 307 370 309
rect 401 307 403 309
rect 418 307 420 309
rect 435 309 437 311
rect 445 309 447 311
rect 468 307 470 309
rect 485 307 487 309
rect 502 309 504 311
rect 512 309 514 311
rect 544 315 546 317
rect 535 302 537 304
rect 554 302 556 304
rect 594 310 596 312
rect 620 315 622 317
rect 606 307 608 309
rect 19 282 21 284
rect 38 282 40 284
rect 28 269 30 271
rect 87 276 89 278
rect 111 277 113 279
rect 97 269 99 271
rect 123 274 125 276
rect 201 276 203 278
rect 225 277 227 279
rect 211 269 213 271
rect 237 274 239 276
rect 282 276 284 278
rect 324 275 326 277
rect 334 275 336 277
rect 351 277 353 279
rect 368 277 370 279
rect 401 277 403 279
rect 418 277 420 279
rect 435 275 437 277
rect 445 275 447 277
rect 468 277 470 279
rect 485 277 487 279
rect 535 282 537 284
rect 502 275 504 277
rect 512 275 514 277
rect 554 282 556 284
rect 544 269 546 271
rect 594 274 596 276
rect 606 277 608 279
rect 620 269 622 271
rect 28 171 30 173
rect 19 158 21 160
rect 97 171 99 173
rect 87 164 89 166
rect 111 163 113 165
rect 38 158 40 160
rect 123 166 125 168
rect 211 171 213 173
rect 201 164 203 166
rect 225 163 227 165
rect 237 166 239 168
rect 282 164 284 166
rect 324 165 326 167
rect 334 165 336 167
rect 351 163 353 165
rect 368 163 370 165
rect 401 163 403 165
rect 418 163 420 165
rect 435 165 437 167
rect 445 165 447 167
rect 468 163 470 165
rect 485 163 487 165
rect 502 165 504 167
rect 512 165 514 167
rect 544 171 546 173
rect 535 158 537 160
rect 554 158 556 160
rect 594 166 596 168
rect 620 171 622 173
rect 606 163 608 165
rect 19 138 21 140
rect 38 138 40 140
rect 28 125 30 127
rect 87 132 89 134
rect 111 133 113 135
rect 97 125 99 127
rect 123 130 125 132
rect 201 132 203 134
rect 225 133 227 135
rect 211 125 213 127
rect 237 130 239 132
rect 282 132 284 134
rect 324 131 326 133
rect 334 131 336 133
rect 351 133 353 135
rect 368 133 370 135
rect 401 133 403 135
rect 418 133 420 135
rect 435 131 437 133
rect 445 131 447 133
rect 468 133 470 135
rect 485 133 487 135
rect 535 138 537 140
rect 502 131 504 133
rect 512 131 514 133
rect 554 138 556 140
rect 544 125 546 127
rect 594 130 596 132
rect 606 133 608 135
rect 620 125 622 127
rect 28 27 30 29
rect 19 14 21 16
rect 97 27 99 29
rect 87 20 89 22
rect 111 19 113 21
rect 38 14 40 16
rect 123 22 125 24
rect 211 27 213 29
rect 201 20 203 22
rect 225 19 227 21
rect 237 22 239 24
rect 282 20 284 22
rect 324 21 326 23
rect 334 21 336 23
rect 351 19 353 21
rect 368 19 370 21
rect 401 19 403 21
rect 418 19 420 21
rect 435 21 437 23
rect 445 21 447 23
rect 468 19 470 21
rect 485 19 487 21
rect 502 21 504 23
rect 512 21 514 23
rect 544 27 546 29
rect 535 14 537 16
rect 554 14 556 16
rect 594 22 596 24
rect 620 27 622 29
rect 606 19 608 21
<< ndifct1 >>
rect 68 574 70 576
rect 8 557 10 559
rect 151 574 153 576
rect 182 574 184 576
rect 57 562 59 564
rect 133 564 135 566
rect 265 574 267 576
rect 301 574 303 576
rect 171 562 173 564
rect 247 564 249 566
rect 312 562 314 564
rect 378 562 380 564
rect 391 562 393 564
rect 458 562 460 564
rect 566 574 568 576
rect 524 557 526 559
rect 584 564 586 566
rect 8 459 10 461
rect 57 454 59 456
rect 133 452 135 454
rect 68 442 70 444
rect 171 454 173 456
rect 151 442 153 444
rect 247 452 249 454
rect 182 442 184 444
rect 312 454 314 456
rect 265 442 267 444
rect 301 442 303 444
rect 378 454 380 456
rect 391 454 393 456
rect 458 454 460 456
rect 524 459 526 461
rect 584 452 586 454
rect 566 442 568 444
rect 68 430 70 432
rect 8 413 10 415
rect 151 430 153 432
rect 182 430 184 432
rect 57 418 59 420
rect 133 420 135 422
rect 265 430 267 432
rect 301 430 303 432
rect 171 418 173 420
rect 247 420 249 422
rect 312 418 314 420
rect 378 418 380 420
rect 391 418 393 420
rect 458 418 460 420
rect 566 430 568 432
rect 524 413 526 415
rect 584 420 586 422
rect 8 315 10 317
rect 57 310 59 312
rect 133 308 135 310
rect 68 298 70 300
rect 171 310 173 312
rect 151 298 153 300
rect 247 308 249 310
rect 182 298 184 300
rect 312 310 314 312
rect 265 298 267 300
rect 301 298 303 300
rect 378 310 380 312
rect 391 310 393 312
rect 458 310 460 312
rect 524 315 526 317
rect 584 308 586 310
rect 566 298 568 300
rect 68 286 70 288
rect 8 269 10 271
rect 151 286 153 288
rect 182 286 184 288
rect 57 274 59 276
rect 133 276 135 278
rect 265 286 267 288
rect 301 286 303 288
rect 171 274 173 276
rect 247 276 249 278
rect 312 274 314 276
rect 378 274 380 276
rect 391 274 393 276
rect 458 274 460 276
rect 566 286 568 288
rect 524 269 526 271
rect 584 276 586 278
rect 8 171 10 173
rect 57 166 59 168
rect 133 164 135 166
rect 68 154 70 156
rect 171 166 173 168
rect 151 154 153 156
rect 247 164 249 166
rect 182 154 184 156
rect 312 166 314 168
rect 265 154 267 156
rect 301 154 303 156
rect 378 166 380 168
rect 391 166 393 168
rect 458 166 460 168
rect 524 171 526 173
rect 584 164 586 166
rect 566 154 568 156
rect 68 142 70 144
rect 8 125 10 127
rect 151 142 153 144
rect 182 142 184 144
rect 57 130 59 132
rect 133 132 135 134
rect 265 142 267 144
rect 301 142 303 144
rect 171 130 173 132
rect 247 132 249 134
rect 312 130 314 132
rect 378 130 380 132
rect 391 130 393 132
rect 458 130 460 132
rect 566 142 568 144
rect 524 125 526 127
rect 584 132 586 134
rect 8 27 10 29
rect 57 22 59 24
rect 133 20 135 22
rect 68 10 70 12
rect 171 22 173 24
rect 151 10 153 12
rect 247 20 249 22
rect 182 10 184 12
rect 312 22 314 24
rect 265 10 267 12
rect 301 10 303 12
rect 378 22 380 24
rect 391 22 393 24
rect 458 22 460 24
rect 524 27 526 29
rect 584 20 586 22
rect 566 10 568 12
<< ntiect1 >>
rect 9 514 11 516
rect 58 514 60 516
rect 131 514 133 516
rect 172 514 174 516
rect 245 514 247 516
rect 311 514 313 516
rect 525 514 527 516
rect 586 514 588 516
rect 9 502 11 504
rect 58 502 60 504
rect 131 502 133 504
rect 172 502 174 504
rect 245 502 247 504
rect 311 502 313 504
rect 525 502 527 504
rect 586 502 588 504
rect 9 370 11 372
rect 58 370 60 372
rect 131 370 133 372
rect 172 370 174 372
rect 245 370 247 372
rect 311 370 313 372
rect 525 370 527 372
rect 586 370 588 372
rect 9 358 11 360
rect 58 358 60 360
rect 131 358 133 360
rect 172 358 174 360
rect 245 358 247 360
rect 311 358 313 360
rect 525 358 527 360
rect 586 358 588 360
rect 9 226 11 228
rect 58 226 60 228
rect 131 226 133 228
rect 172 226 174 228
rect 245 226 247 228
rect 311 226 313 228
rect 525 226 527 228
rect 586 226 588 228
rect 9 214 11 216
rect 58 214 60 216
rect 131 214 133 216
rect 172 214 174 216
rect 245 214 247 216
rect 311 214 313 216
rect 525 214 527 216
rect 586 214 588 216
rect 9 82 11 84
rect 58 82 60 84
rect 131 82 133 84
rect 172 82 174 84
rect 245 82 247 84
rect 311 82 313 84
rect 525 82 527 84
rect 586 82 588 84
rect 9 70 11 72
rect 58 70 60 72
rect 131 70 133 72
rect 172 70 174 72
rect 245 70 247 72
rect 311 70 313 72
rect 525 70 527 72
rect 586 70 588 72
<< ptiect1 >>
rect 9 574 11 576
rect 58 574 60 576
rect 98 574 100 576
rect 172 574 174 576
rect 212 574 214 576
rect 311 574 313 576
rect 525 574 527 576
rect 619 574 621 576
rect 9 442 11 444
rect 58 442 60 444
rect 98 442 100 444
rect 172 442 174 444
rect 212 442 214 444
rect 311 442 313 444
rect 525 442 527 444
rect 619 442 621 444
rect 9 430 11 432
rect 58 430 60 432
rect 98 430 100 432
rect 172 430 174 432
rect 212 430 214 432
rect 311 430 313 432
rect 525 430 527 432
rect 619 430 621 432
rect 9 298 11 300
rect 58 298 60 300
rect 98 298 100 300
rect 172 298 174 300
rect 212 298 214 300
rect 311 298 313 300
rect 525 298 527 300
rect 619 298 621 300
rect 9 286 11 288
rect 58 286 60 288
rect 98 286 100 288
rect 172 286 174 288
rect 212 286 214 288
rect 311 286 313 288
rect 525 286 527 288
rect 619 286 621 288
rect 9 154 11 156
rect 58 154 60 156
rect 98 154 100 156
rect 172 154 174 156
rect 212 154 214 156
rect 311 154 313 156
rect 525 154 527 156
rect 619 154 621 156
rect 9 142 11 144
rect 58 142 60 144
rect 98 142 100 144
rect 172 142 174 144
rect 212 142 214 144
rect 311 142 313 144
rect 525 142 527 144
rect 619 142 621 144
rect 9 10 11 12
rect 58 10 60 12
rect 98 10 100 12
rect 172 10 174 12
rect 212 10 214 12
rect 311 10 313 12
rect 525 10 527 12
rect 619 10 621 12
<< pdifct0 >>
rect 19 517 21 519
rect 38 524 40 526
rect 105 538 107 540
rect 67 526 69 528
rect 77 531 79 533
rect 77 524 79 526
rect 87 524 89 526
rect 115 524 117 526
rect 131 538 133 540
rect 131 531 133 533
rect 115 517 117 519
rect 151 523 153 525
rect 219 538 221 540
rect 181 526 183 528
rect 191 531 193 533
rect 191 524 193 526
rect 201 524 203 526
rect 229 524 231 526
rect 245 538 247 540
rect 245 531 247 533
rect 229 517 231 519
rect 265 523 267 525
rect 282 524 284 526
rect 292 531 294 533
rect 292 524 294 526
rect 302 526 304 528
rect 324 539 326 541
rect 334 517 336 519
rect 351 527 353 529
rect 368 517 370 519
rect 445 539 447 541
rect 401 517 403 519
rect 418 527 420 529
rect 435 517 437 519
rect 512 539 514 541
rect 468 517 470 519
rect 485 527 487 529
rect 502 517 504 519
rect 535 517 537 519
rect 554 524 556 526
rect 566 523 568 525
rect 586 538 588 540
rect 586 531 588 533
rect 602 524 604 526
rect 602 517 604 519
rect 612 538 614 540
rect 19 499 21 501
rect 38 492 40 494
rect 67 490 69 492
rect 77 492 79 494
rect 77 485 79 487
rect 87 492 89 494
rect 105 478 107 480
rect 115 499 117 501
rect 115 492 117 494
rect 131 485 133 487
rect 131 478 133 480
rect 151 493 153 495
rect 181 490 183 492
rect 191 492 193 494
rect 191 485 193 487
rect 201 492 203 494
rect 219 478 221 480
rect 229 499 231 501
rect 229 492 231 494
rect 245 485 247 487
rect 245 478 247 480
rect 334 499 336 501
rect 265 493 267 495
rect 282 492 284 494
rect 292 492 294 494
rect 292 485 294 487
rect 302 490 304 492
rect 351 489 353 491
rect 368 499 370 501
rect 324 477 326 479
rect 401 499 403 501
rect 418 489 420 491
rect 435 499 437 501
rect 468 499 470 501
rect 485 489 487 491
rect 502 499 504 501
rect 535 499 537 501
rect 445 477 447 479
rect 512 477 514 479
rect 554 492 556 494
rect 566 493 568 495
rect 602 499 604 501
rect 586 485 588 487
rect 586 478 588 480
rect 602 492 604 494
rect 612 478 614 480
rect 19 373 21 375
rect 38 380 40 382
rect 105 394 107 396
rect 67 382 69 384
rect 77 387 79 389
rect 77 380 79 382
rect 87 380 89 382
rect 115 380 117 382
rect 131 394 133 396
rect 131 387 133 389
rect 115 373 117 375
rect 151 379 153 381
rect 219 394 221 396
rect 181 382 183 384
rect 191 387 193 389
rect 191 380 193 382
rect 201 380 203 382
rect 229 380 231 382
rect 245 394 247 396
rect 245 387 247 389
rect 229 373 231 375
rect 265 379 267 381
rect 282 380 284 382
rect 292 387 294 389
rect 292 380 294 382
rect 302 382 304 384
rect 324 395 326 397
rect 334 373 336 375
rect 351 383 353 385
rect 368 373 370 375
rect 445 395 447 397
rect 401 373 403 375
rect 418 383 420 385
rect 435 373 437 375
rect 512 395 514 397
rect 468 373 470 375
rect 485 383 487 385
rect 502 373 504 375
rect 535 373 537 375
rect 554 380 556 382
rect 566 379 568 381
rect 586 394 588 396
rect 586 387 588 389
rect 602 380 604 382
rect 602 373 604 375
rect 612 394 614 396
rect 19 355 21 357
rect 38 348 40 350
rect 67 346 69 348
rect 77 348 79 350
rect 77 341 79 343
rect 87 348 89 350
rect 105 334 107 336
rect 115 355 117 357
rect 115 348 117 350
rect 131 341 133 343
rect 131 334 133 336
rect 151 349 153 351
rect 181 346 183 348
rect 191 348 193 350
rect 191 341 193 343
rect 201 348 203 350
rect 219 334 221 336
rect 229 355 231 357
rect 229 348 231 350
rect 245 341 247 343
rect 245 334 247 336
rect 334 355 336 357
rect 265 349 267 351
rect 282 348 284 350
rect 292 348 294 350
rect 292 341 294 343
rect 302 346 304 348
rect 351 345 353 347
rect 368 355 370 357
rect 324 333 326 335
rect 401 355 403 357
rect 418 345 420 347
rect 435 355 437 357
rect 468 355 470 357
rect 485 345 487 347
rect 502 355 504 357
rect 535 355 537 357
rect 445 333 447 335
rect 512 333 514 335
rect 554 348 556 350
rect 566 349 568 351
rect 602 355 604 357
rect 586 341 588 343
rect 586 334 588 336
rect 602 348 604 350
rect 612 334 614 336
rect 19 229 21 231
rect 38 236 40 238
rect 105 250 107 252
rect 67 238 69 240
rect 77 243 79 245
rect 77 236 79 238
rect 87 236 89 238
rect 115 236 117 238
rect 131 250 133 252
rect 131 243 133 245
rect 115 229 117 231
rect 151 235 153 237
rect 219 250 221 252
rect 181 238 183 240
rect 191 243 193 245
rect 191 236 193 238
rect 201 236 203 238
rect 229 236 231 238
rect 245 250 247 252
rect 245 243 247 245
rect 229 229 231 231
rect 265 235 267 237
rect 282 236 284 238
rect 292 243 294 245
rect 292 236 294 238
rect 302 238 304 240
rect 324 251 326 253
rect 334 229 336 231
rect 351 239 353 241
rect 368 229 370 231
rect 445 251 447 253
rect 401 229 403 231
rect 418 239 420 241
rect 435 229 437 231
rect 512 251 514 253
rect 468 229 470 231
rect 485 239 487 241
rect 502 229 504 231
rect 535 229 537 231
rect 554 236 556 238
rect 566 235 568 237
rect 586 250 588 252
rect 586 243 588 245
rect 602 236 604 238
rect 602 229 604 231
rect 612 250 614 252
rect 19 211 21 213
rect 38 204 40 206
rect 67 202 69 204
rect 77 204 79 206
rect 77 197 79 199
rect 87 204 89 206
rect 105 190 107 192
rect 115 211 117 213
rect 115 204 117 206
rect 131 197 133 199
rect 131 190 133 192
rect 151 205 153 207
rect 181 202 183 204
rect 191 204 193 206
rect 191 197 193 199
rect 201 204 203 206
rect 219 190 221 192
rect 229 211 231 213
rect 229 204 231 206
rect 245 197 247 199
rect 245 190 247 192
rect 334 211 336 213
rect 265 205 267 207
rect 282 204 284 206
rect 292 204 294 206
rect 292 197 294 199
rect 302 202 304 204
rect 351 201 353 203
rect 368 211 370 213
rect 324 189 326 191
rect 401 211 403 213
rect 418 201 420 203
rect 435 211 437 213
rect 468 211 470 213
rect 485 201 487 203
rect 502 211 504 213
rect 535 211 537 213
rect 445 189 447 191
rect 512 189 514 191
rect 554 204 556 206
rect 566 205 568 207
rect 602 211 604 213
rect 586 197 588 199
rect 586 190 588 192
rect 602 204 604 206
rect 612 190 614 192
rect 19 85 21 87
rect 38 92 40 94
rect 105 106 107 108
rect 67 94 69 96
rect 77 99 79 101
rect 77 92 79 94
rect 87 92 89 94
rect 115 92 117 94
rect 131 106 133 108
rect 131 99 133 101
rect 115 85 117 87
rect 151 91 153 93
rect 219 106 221 108
rect 181 94 183 96
rect 191 99 193 101
rect 191 92 193 94
rect 201 92 203 94
rect 229 92 231 94
rect 245 106 247 108
rect 245 99 247 101
rect 229 85 231 87
rect 265 91 267 93
rect 282 92 284 94
rect 292 99 294 101
rect 292 92 294 94
rect 302 94 304 96
rect 324 107 326 109
rect 334 85 336 87
rect 351 95 353 97
rect 368 85 370 87
rect 445 107 447 109
rect 401 85 403 87
rect 418 95 420 97
rect 435 85 437 87
rect 512 107 514 109
rect 468 85 470 87
rect 485 95 487 97
rect 502 85 504 87
rect 535 85 537 87
rect 554 92 556 94
rect 566 91 568 93
rect 586 106 588 108
rect 586 99 588 101
rect 602 92 604 94
rect 602 85 604 87
rect 612 106 614 108
rect 19 67 21 69
rect 38 60 40 62
rect 67 58 69 60
rect 77 60 79 62
rect 77 53 79 55
rect 87 60 89 62
rect 105 46 107 48
rect 115 67 117 69
rect 115 60 117 62
rect 131 53 133 55
rect 131 46 133 48
rect 151 61 153 63
rect 181 58 183 60
rect 191 60 193 62
rect 191 53 193 55
rect 201 60 203 62
rect 219 46 221 48
rect 229 67 231 69
rect 229 60 231 62
rect 245 53 247 55
rect 245 46 247 48
rect 334 67 336 69
rect 265 61 267 63
rect 282 60 284 62
rect 292 60 294 62
rect 292 53 294 55
rect 302 58 304 60
rect 351 57 353 59
rect 368 67 370 69
rect 324 45 326 47
rect 401 67 403 69
rect 418 57 420 59
rect 435 67 437 69
rect 468 67 470 69
rect 485 57 487 59
rect 502 67 504 69
rect 535 67 537 69
rect 445 45 447 47
rect 512 45 514 47
rect 554 60 556 62
rect 566 61 568 63
rect 602 67 604 69
rect 586 53 588 55
rect 586 46 588 48
rect 602 60 604 62
rect 612 46 614 48
<< pdifct1 >>
rect 8 534 10 536
rect 8 527 10 529
rect 57 538 59 540
rect 57 531 59 533
rect 141 531 143 533
rect 171 538 173 540
rect 171 531 173 533
rect 255 531 257 533
rect 312 538 314 540
rect 312 531 314 533
rect 378 524 380 526
rect 391 524 393 526
rect 458 524 460 526
rect 524 534 526 536
rect 524 527 526 529
rect 576 531 578 533
rect 8 489 10 491
rect 8 482 10 484
rect 57 485 59 487
rect 57 478 59 480
rect 141 485 143 487
rect 171 485 173 487
rect 171 478 173 480
rect 255 485 257 487
rect 312 485 314 487
rect 312 478 314 480
rect 378 492 380 494
rect 391 492 393 494
rect 458 492 460 494
rect 524 489 526 491
rect 524 482 526 484
rect 576 485 578 487
rect 8 390 10 392
rect 8 383 10 385
rect 57 394 59 396
rect 57 387 59 389
rect 141 387 143 389
rect 171 394 173 396
rect 171 387 173 389
rect 255 387 257 389
rect 312 394 314 396
rect 312 387 314 389
rect 378 380 380 382
rect 391 380 393 382
rect 458 380 460 382
rect 524 390 526 392
rect 524 383 526 385
rect 576 387 578 389
rect 8 345 10 347
rect 8 338 10 340
rect 57 341 59 343
rect 57 334 59 336
rect 141 341 143 343
rect 171 341 173 343
rect 171 334 173 336
rect 255 341 257 343
rect 312 341 314 343
rect 312 334 314 336
rect 378 348 380 350
rect 391 348 393 350
rect 458 348 460 350
rect 524 345 526 347
rect 524 338 526 340
rect 576 341 578 343
rect 8 246 10 248
rect 8 239 10 241
rect 57 250 59 252
rect 57 243 59 245
rect 141 243 143 245
rect 171 250 173 252
rect 171 243 173 245
rect 255 243 257 245
rect 312 250 314 252
rect 312 243 314 245
rect 378 236 380 238
rect 391 236 393 238
rect 458 236 460 238
rect 524 246 526 248
rect 524 239 526 241
rect 576 243 578 245
rect 8 201 10 203
rect 8 194 10 196
rect 57 197 59 199
rect 57 190 59 192
rect 141 197 143 199
rect 171 197 173 199
rect 171 190 173 192
rect 255 197 257 199
rect 312 197 314 199
rect 312 190 314 192
rect 378 204 380 206
rect 391 204 393 206
rect 458 204 460 206
rect 524 201 526 203
rect 524 194 526 196
rect 576 197 578 199
rect 8 102 10 104
rect 8 95 10 97
rect 57 106 59 108
rect 57 99 59 101
rect 141 99 143 101
rect 171 106 173 108
rect 171 99 173 101
rect 255 99 257 101
rect 312 106 314 108
rect 312 99 314 101
rect 378 92 380 94
rect 391 92 393 94
rect 458 92 460 94
rect 524 102 526 104
rect 524 95 526 97
rect 576 99 578 101
rect 8 57 10 59
rect 8 50 10 52
rect 57 53 59 55
rect 57 46 59 48
rect 141 53 143 55
rect 171 53 173 55
rect 171 46 173 48
rect 255 53 257 55
rect 312 53 314 55
rect 312 46 314 48
rect 378 60 380 62
rect 391 60 393 62
rect 458 60 460 62
rect 524 57 526 59
rect 524 50 526 52
rect 576 53 578 55
<< alu0 >>
rect 17 572 23 573
rect 17 570 19 572
rect 21 570 23 572
rect 17 569 23 570
rect 36 572 42 573
rect 36 570 38 572
rect 40 570 42 572
rect 36 569 42 570
rect 109 567 115 573
rect 71 566 91 567
rect 71 564 87 566
rect 89 564 91 566
rect 109 565 111 567
rect 113 565 115 567
rect 109 564 115 565
rect 122 564 126 566
rect 71 563 91 564
rect 14 559 32 560
rect 14 557 28 559
rect 30 557 32 559
rect 14 556 32 557
rect 14 550 18 556
rect 14 548 15 550
rect 17 548 18 550
rect 10 527 11 538
rect 14 535 18 548
rect 33 543 39 544
rect 59 560 60 562
rect 71 559 75 563
rect 122 562 123 564
rect 125 562 126 564
rect 63 555 75 559
rect 63 550 67 555
rect 63 548 64 550
rect 66 548 67 550
rect 14 531 29 535
rect 25 527 29 531
rect 63 536 67 548
rect 96 559 100 561
rect 96 557 97 559
rect 99 557 100 559
rect 96 551 100 557
rect 122 559 126 562
rect 122 555 146 559
rect 96 547 107 551
rect 63 533 80 536
rect 63 532 77 533
rect 76 531 77 532
rect 79 531 80 533
rect 65 528 71 529
rect 25 526 42 527
rect 25 524 38 526
rect 40 524 42 526
rect 25 523 42 524
rect 65 526 67 528
rect 69 526 71 528
rect 17 519 23 520
rect 17 517 19 519
rect 21 517 23 519
rect 65 517 71 526
rect 76 526 80 531
rect 103 541 107 547
rect 142 551 146 555
rect 122 550 138 551
rect 122 548 134 550
rect 136 548 138 550
rect 122 547 138 548
rect 142 549 147 551
rect 142 547 144 549
rect 146 547 147 549
rect 122 541 126 547
rect 142 545 147 547
rect 142 543 146 545
rect 103 540 126 541
rect 103 538 105 540
rect 107 538 126 540
rect 103 537 126 538
rect 76 524 77 526
rect 79 524 80 526
rect 76 522 80 524
rect 85 526 91 527
rect 85 524 87 526
rect 89 524 91 526
rect 85 517 91 524
rect 114 526 118 528
rect 114 524 115 526
rect 117 524 118 526
rect 114 519 118 524
rect 122 526 126 537
rect 130 540 146 543
rect 130 538 131 540
rect 133 539 146 540
rect 133 538 134 539
rect 130 533 134 538
rect 130 531 131 533
rect 133 531 134 533
rect 130 529 134 531
rect 223 567 229 573
rect 185 566 205 567
rect 185 564 201 566
rect 203 564 205 566
rect 223 565 225 567
rect 227 565 229 567
rect 223 564 229 565
rect 236 564 240 566
rect 185 563 205 564
rect 173 560 174 562
rect 185 559 189 563
rect 236 562 237 564
rect 239 562 240 564
rect 280 566 300 567
rect 280 564 282 566
rect 284 564 300 566
rect 280 563 300 564
rect 177 555 189 559
rect 177 550 181 555
rect 177 548 178 550
rect 180 548 181 550
rect 177 536 181 548
rect 210 559 214 561
rect 210 557 211 559
rect 213 557 214 559
rect 210 551 214 557
rect 236 559 240 562
rect 236 555 260 559
rect 210 547 221 551
rect 177 533 194 536
rect 177 532 191 533
rect 190 531 191 532
rect 193 531 194 533
rect 179 528 185 529
rect 179 526 181 528
rect 183 526 185 528
rect 122 525 155 526
rect 122 523 151 525
rect 153 523 155 525
rect 122 522 155 523
rect 114 517 115 519
rect 117 517 118 519
rect 179 517 185 526
rect 190 526 194 531
rect 217 541 221 547
rect 256 551 260 555
rect 236 550 252 551
rect 236 548 248 550
rect 250 548 252 550
rect 236 547 252 548
rect 256 549 261 551
rect 256 547 258 549
rect 260 547 261 549
rect 236 541 240 547
rect 256 545 261 547
rect 256 543 260 545
rect 217 540 240 541
rect 217 538 219 540
rect 221 538 240 540
rect 217 537 240 538
rect 190 524 191 526
rect 193 524 194 526
rect 190 522 194 524
rect 199 526 205 527
rect 199 524 201 526
rect 203 524 205 526
rect 199 517 205 524
rect 228 526 232 528
rect 228 524 229 526
rect 231 524 232 526
rect 228 519 232 524
rect 236 526 240 537
rect 244 540 260 543
rect 244 538 245 540
rect 247 539 260 540
rect 296 559 300 563
rect 311 560 312 562
rect 296 555 308 559
rect 304 550 308 555
rect 304 548 305 550
rect 307 548 308 550
rect 247 538 248 539
rect 244 533 248 538
rect 244 531 245 533
rect 247 531 248 533
rect 244 529 248 531
rect 304 536 308 548
rect 291 533 308 536
rect 291 531 292 533
rect 294 532 308 533
rect 322 565 328 566
rect 322 563 324 565
rect 326 563 328 565
rect 322 562 328 563
rect 332 565 338 573
rect 332 563 334 565
rect 336 563 338 565
rect 349 567 364 568
rect 349 565 351 567
rect 353 565 364 567
rect 349 564 364 565
rect 332 562 338 563
rect 322 542 326 562
rect 360 559 364 564
rect 367 567 371 573
rect 367 565 368 567
rect 370 565 371 567
rect 367 563 371 565
rect 346 556 357 558
rect 346 554 354 556
rect 356 554 357 556
rect 360 557 374 559
rect 360 555 375 557
rect 346 552 357 554
rect 370 553 372 555
rect 374 553 375 555
rect 346 542 350 552
rect 370 551 375 553
rect 322 541 350 542
rect 322 539 324 541
rect 326 540 350 541
rect 326 539 347 540
rect 322 538 347 539
rect 349 538 350 540
rect 366 541 367 547
rect 346 536 350 538
rect 294 531 295 532
rect 280 526 286 527
rect 236 525 269 526
rect 236 523 265 525
rect 267 523 269 525
rect 236 522 269 523
rect 280 524 282 526
rect 284 524 286 526
rect 228 517 229 519
rect 231 517 232 519
rect 280 517 286 524
rect 291 526 295 531
rect 370 534 374 551
rect 358 530 374 534
rect 291 524 292 526
rect 294 524 295 526
rect 291 522 295 524
rect 300 528 306 529
rect 300 526 302 528
rect 304 526 306 528
rect 300 517 306 526
rect 349 529 362 530
rect 349 527 351 529
rect 353 527 362 529
rect 349 526 362 527
rect 400 567 404 573
rect 400 565 401 567
rect 403 565 404 567
rect 400 563 404 565
rect 407 567 422 568
rect 407 565 418 567
rect 420 565 422 567
rect 407 564 422 565
rect 433 565 439 573
rect 467 567 471 573
rect 407 559 411 564
rect 433 563 435 565
rect 437 563 439 565
rect 433 562 439 563
rect 443 565 449 566
rect 443 563 445 565
rect 447 563 449 565
rect 443 562 449 563
rect 397 557 411 559
rect 396 555 411 557
rect 414 556 425 558
rect 396 553 397 555
rect 399 553 401 555
rect 396 551 401 553
rect 414 554 415 556
rect 417 554 425 556
rect 414 552 425 554
rect 397 534 401 551
rect 404 541 405 547
rect 421 542 425 552
rect 445 542 449 562
rect 421 541 449 542
rect 421 540 445 541
rect 421 538 422 540
rect 424 539 445 540
rect 447 539 449 541
rect 424 538 449 539
rect 467 565 468 567
rect 470 565 471 567
rect 467 563 471 565
rect 474 567 489 568
rect 474 565 485 567
rect 487 565 489 567
rect 474 564 489 565
rect 500 565 506 573
rect 533 572 539 573
rect 533 570 535 572
rect 537 570 539 572
rect 533 569 539 570
rect 552 572 558 573
rect 552 570 554 572
rect 556 570 558 572
rect 552 569 558 570
rect 604 567 610 573
rect 474 559 478 564
rect 500 563 502 565
rect 504 563 506 565
rect 500 562 506 563
rect 510 565 516 566
rect 510 563 512 565
rect 514 563 516 565
rect 510 562 516 563
rect 464 557 478 559
rect 421 536 425 538
rect 397 530 413 534
rect 409 529 422 530
rect 409 527 418 529
rect 420 527 422 529
rect 409 526 422 527
rect 463 555 478 557
rect 481 556 492 558
rect 463 553 464 555
rect 466 553 468 555
rect 463 551 468 553
rect 481 554 482 556
rect 484 554 492 556
rect 481 552 492 554
rect 464 534 468 551
rect 471 541 472 547
rect 488 542 492 552
rect 512 542 516 562
rect 593 564 597 566
rect 604 565 606 567
rect 608 565 610 567
rect 604 564 610 565
rect 488 541 516 542
rect 488 540 512 541
rect 488 538 489 540
rect 491 539 512 540
rect 514 539 516 541
rect 491 538 516 539
rect 530 559 548 560
rect 530 557 544 559
rect 546 557 548 559
rect 530 556 548 557
rect 488 536 492 538
rect 530 550 534 556
rect 530 548 531 550
rect 533 548 534 550
rect 464 530 480 534
rect 476 529 489 530
rect 476 527 485 529
rect 487 527 489 529
rect 476 526 489 527
rect 526 527 527 538
rect 530 535 534 548
rect 593 562 594 564
rect 596 562 597 564
rect 593 559 597 562
rect 549 543 555 544
rect 530 531 545 535
rect 541 527 545 531
rect 573 555 597 559
rect 573 551 577 555
rect 619 559 623 561
rect 619 557 620 559
rect 622 557 623 559
rect 572 549 577 551
rect 572 547 573 549
rect 575 547 577 549
rect 581 550 597 551
rect 581 548 583 550
rect 585 548 597 550
rect 581 547 597 548
rect 572 545 577 547
rect 573 543 577 545
rect 573 540 589 543
rect 573 539 586 540
rect 585 538 586 539
rect 588 538 589 540
rect 585 533 589 538
rect 585 531 586 533
rect 588 531 589 533
rect 585 529 589 531
rect 593 541 597 547
rect 619 551 623 557
rect 612 547 623 551
rect 612 541 616 547
rect 593 540 616 541
rect 593 538 612 540
rect 614 538 616 540
rect 593 537 616 538
rect 541 526 558 527
rect 593 526 597 537
rect 541 524 554 526
rect 556 524 558 526
rect 541 523 558 524
rect 564 525 597 526
rect 564 523 566 525
rect 568 523 597 525
rect 564 522 597 523
rect 601 526 605 528
rect 601 524 602 526
rect 604 524 605 526
rect 333 519 337 521
rect 333 517 334 519
rect 336 517 337 519
rect 366 519 372 520
rect 366 517 368 519
rect 370 517 372 519
rect 399 519 405 520
rect 399 517 401 519
rect 403 517 405 519
rect 434 519 438 521
rect 434 517 435 519
rect 437 517 438 519
rect 466 519 472 520
rect 466 517 468 519
rect 470 517 472 519
rect 501 519 505 521
rect 501 517 502 519
rect 504 517 505 519
rect 533 519 539 520
rect 533 517 535 519
rect 537 517 539 519
rect 601 519 605 524
rect 601 517 602 519
rect 604 517 605 519
rect 17 499 19 501
rect 21 499 23 501
rect 17 498 23 499
rect 25 494 42 495
rect 25 492 38 494
rect 40 492 42 494
rect 25 491 42 492
rect 65 492 71 501
rect 10 480 11 491
rect 25 487 29 491
rect 65 490 67 492
rect 69 490 71 492
rect 65 489 71 490
rect 76 494 80 496
rect 76 492 77 494
rect 79 492 80 494
rect 14 483 29 487
rect 76 487 80 492
rect 85 494 91 501
rect 114 499 115 501
rect 117 499 118 501
rect 85 492 87 494
rect 89 492 91 494
rect 85 491 91 492
rect 114 494 118 499
rect 114 492 115 494
rect 117 492 118 494
rect 114 490 118 492
rect 122 495 155 496
rect 122 493 151 495
rect 153 493 155 495
rect 122 492 155 493
rect 179 492 185 501
rect 76 486 77 487
rect 14 470 18 483
rect 63 485 77 486
rect 79 485 80 487
rect 63 482 80 485
rect 33 474 39 475
rect 14 468 15 470
rect 17 468 18 470
rect 14 462 18 468
rect 14 461 32 462
rect 14 459 28 461
rect 30 459 32 461
rect 14 458 32 459
rect 63 470 67 482
rect 122 481 126 492
rect 179 490 181 492
rect 183 490 185 492
rect 179 489 185 490
rect 190 494 194 496
rect 190 492 191 494
rect 193 492 194 494
rect 103 480 126 481
rect 103 478 105 480
rect 107 478 126 480
rect 103 477 126 478
rect 103 471 107 477
rect 63 468 64 470
rect 66 468 67 470
rect 63 463 67 468
rect 63 459 75 463
rect 59 456 60 458
rect 71 455 75 459
rect 96 467 107 471
rect 96 461 100 467
rect 122 471 126 477
rect 130 487 134 489
rect 130 485 131 487
rect 133 485 134 487
rect 130 480 134 485
rect 130 478 131 480
rect 133 479 134 480
rect 133 478 146 479
rect 130 475 146 478
rect 142 473 146 475
rect 142 471 147 473
rect 122 470 138 471
rect 122 468 134 470
rect 136 468 138 470
rect 122 467 138 468
rect 142 469 144 471
rect 146 469 147 471
rect 142 467 147 469
rect 96 459 97 461
rect 99 459 100 461
rect 96 457 100 459
rect 142 463 146 467
rect 122 459 146 463
rect 122 456 126 459
rect 71 454 91 455
rect 122 454 123 456
rect 125 454 126 456
rect 71 452 87 454
rect 89 452 91 454
rect 71 451 91 452
rect 109 453 115 454
rect 109 451 111 453
rect 113 451 115 453
rect 122 452 126 454
rect 190 487 194 492
rect 199 494 205 501
rect 228 499 229 501
rect 231 499 232 501
rect 199 492 201 494
rect 203 492 205 494
rect 199 491 205 492
rect 228 494 232 499
rect 228 492 229 494
rect 231 492 232 494
rect 228 490 232 492
rect 236 495 269 496
rect 236 493 265 495
rect 267 493 269 495
rect 236 492 269 493
rect 280 494 286 501
rect 280 492 282 494
rect 284 492 286 494
rect 190 486 191 487
rect 177 485 191 486
rect 193 485 194 487
rect 177 482 194 485
rect 177 470 181 482
rect 236 481 240 492
rect 280 491 286 492
rect 291 494 295 496
rect 291 492 292 494
rect 294 492 295 494
rect 217 480 240 481
rect 217 478 219 480
rect 221 478 240 480
rect 217 477 240 478
rect 217 471 221 477
rect 177 468 178 470
rect 180 468 181 470
rect 177 463 181 468
rect 177 459 189 463
rect 173 456 174 458
rect 17 448 23 449
rect 17 446 19 448
rect 21 446 23 448
rect 17 445 23 446
rect 36 448 42 449
rect 36 446 38 448
rect 40 446 42 448
rect 36 445 42 446
rect 109 445 115 451
rect 185 455 189 459
rect 210 467 221 471
rect 210 461 214 467
rect 236 471 240 477
rect 244 487 248 489
rect 244 485 245 487
rect 247 485 248 487
rect 244 480 248 485
rect 244 478 245 480
rect 247 479 248 480
rect 247 478 260 479
rect 244 475 260 478
rect 256 473 260 475
rect 291 487 295 492
rect 300 492 306 501
rect 333 499 334 501
rect 336 499 337 501
rect 333 497 337 499
rect 366 499 368 501
rect 370 499 372 501
rect 366 498 372 499
rect 399 499 401 501
rect 403 499 405 501
rect 399 498 405 499
rect 434 499 435 501
rect 437 499 438 501
rect 434 497 438 499
rect 466 499 468 501
rect 470 499 472 501
rect 466 498 472 499
rect 501 499 502 501
rect 504 499 505 501
rect 501 497 505 499
rect 533 499 535 501
rect 537 499 539 501
rect 533 498 539 499
rect 601 499 602 501
rect 604 499 605 501
rect 300 490 302 492
rect 304 490 306 492
rect 300 489 306 490
rect 291 485 292 487
rect 294 486 295 487
rect 294 485 308 486
rect 291 482 308 485
rect 256 471 261 473
rect 236 470 252 471
rect 236 468 248 470
rect 250 468 252 470
rect 236 467 252 468
rect 256 469 258 471
rect 260 469 261 471
rect 256 467 261 469
rect 210 459 211 461
rect 213 459 214 461
rect 210 457 214 459
rect 256 463 260 467
rect 236 459 260 463
rect 236 456 240 459
rect 185 454 205 455
rect 236 454 237 456
rect 239 454 240 456
rect 304 470 308 482
rect 349 491 362 492
rect 349 489 351 491
rect 353 489 362 491
rect 349 488 362 489
rect 358 484 374 488
rect 346 480 350 482
rect 304 468 305 470
rect 307 468 308 470
rect 304 463 308 468
rect 296 459 308 463
rect 296 455 300 459
rect 311 456 312 458
rect 185 452 201 454
rect 203 452 205 454
rect 185 451 205 452
rect 223 453 229 454
rect 223 451 225 453
rect 227 451 229 453
rect 236 452 240 454
rect 280 454 300 455
rect 280 452 282 454
rect 284 452 300 454
rect 280 451 300 452
rect 223 445 229 451
rect 322 479 347 480
rect 322 477 324 479
rect 326 478 347 479
rect 349 478 350 480
rect 326 477 350 478
rect 322 476 350 477
rect 322 456 326 476
rect 346 466 350 476
rect 366 471 367 477
rect 370 467 374 484
rect 346 464 357 466
rect 346 462 354 464
rect 356 462 357 464
rect 370 465 375 467
rect 370 463 372 465
rect 374 463 375 465
rect 346 460 357 462
rect 360 461 375 463
rect 360 459 374 461
rect 322 455 328 456
rect 322 453 324 455
rect 326 453 328 455
rect 322 452 328 453
rect 332 455 338 456
rect 332 453 334 455
rect 336 453 338 455
rect 360 454 364 459
rect 332 445 338 453
rect 349 453 364 454
rect 349 451 351 453
rect 353 451 364 453
rect 349 450 364 451
rect 367 453 371 455
rect 367 451 368 453
rect 370 451 371 453
rect 367 445 371 451
rect 409 491 422 492
rect 409 489 418 491
rect 420 489 422 491
rect 409 488 422 489
rect 397 484 413 488
rect 397 467 401 484
rect 476 491 489 492
rect 421 480 425 482
rect 404 471 405 477
rect 421 478 422 480
rect 424 479 449 480
rect 424 478 445 479
rect 421 477 445 478
rect 447 477 449 479
rect 421 476 449 477
rect 396 465 401 467
rect 421 466 425 476
rect 396 463 397 465
rect 399 463 401 465
rect 414 464 425 466
rect 396 461 411 463
rect 397 459 411 461
rect 414 462 415 464
rect 417 462 425 464
rect 414 460 425 462
rect 400 453 404 455
rect 400 451 401 453
rect 403 451 404 453
rect 400 445 404 451
rect 407 454 411 459
rect 445 456 449 476
rect 433 455 439 456
rect 407 453 422 454
rect 407 451 418 453
rect 420 451 422 453
rect 407 450 422 451
rect 433 453 435 455
rect 437 453 439 455
rect 433 445 439 453
rect 443 455 449 456
rect 443 453 445 455
rect 447 453 449 455
rect 443 452 449 453
rect 476 489 485 491
rect 487 489 489 491
rect 476 488 489 489
rect 464 484 480 488
rect 464 467 468 484
rect 564 495 597 496
rect 541 494 558 495
rect 541 492 554 494
rect 556 492 558 494
rect 564 493 566 495
rect 568 493 597 495
rect 564 492 597 493
rect 541 491 558 492
rect 488 480 492 482
rect 471 471 472 477
rect 488 478 489 480
rect 491 479 516 480
rect 491 478 512 479
rect 488 477 512 478
rect 514 477 516 479
rect 488 476 516 477
rect 463 465 468 467
rect 488 466 492 476
rect 463 463 464 465
rect 466 463 468 465
rect 481 464 492 466
rect 463 461 478 463
rect 464 459 478 461
rect 481 462 482 464
rect 484 462 492 464
rect 481 460 492 462
rect 467 453 471 455
rect 467 451 468 453
rect 470 451 471 453
rect 467 445 471 451
rect 474 454 478 459
rect 512 456 516 476
rect 526 480 527 491
rect 541 487 545 491
rect 530 483 545 487
rect 530 470 534 483
rect 585 487 589 489
rect 585 485 586 487
rect 588 485 589 487
rect 549 474 555 475
rect 530 468 531 470
rect 533 468 534 470
rect 530 462 534 468
rect 530 461 548 462
rect 530 459 544 461
rect 546 459 548 461
rect 530 458 548 459
rect 585 480 589 485
rect 585 479 586 480
rect 573 478 586 479
rect 588 478 589 480
rect 573 475 589 478
rect 593 481 597 492
rect 601 494 605 499
rect 601 492 602 494
rect 604 492 605 494
rect 601 490 605 492
rect 593 480 616 481
rect 593 478 612 480
rect 614 478 616 480
rect 593 477 616 478
rect 573 473 577 475
rect 572 471 577 473
rect 593 471 597 477
rect 572 469 573 471
rect 575 469 577 471
rect 572 467 577 469
rect 581 470 597 471
rect 581 468 583 470
rect 585 468 597 470
rect 581 467 597 468
rect 500 455 506 456
rect 474 453 489 454
rect 474 451 485 453
rect 487 451 489 453
rect 474 450 489 451
rect 500 453 502 455
rect 504 453 506 455
rect 500 445 506 453
rect 510 455 516 456
rect 510 453 512 455
rect 514 453 516 455
rect 510 452 516 453
rect 573 463 577 467
rect 612 471 616 477
rect 612 467 623 471
rect 573 459 597 463
rect 593 456 597 459
rect 619 461 623 467
rect 619 459 620 461
rect 622 459 623 461
rect 619 457 623 459
rect 593 454 594 456
rect 596 454 597 456
rect 593 452 597 454
rect 604 453 610 454
rect 604 451 606 453
rect 608 451 610 453
rect 533 448 539 449
rect 533 446 535 448
rect 537 446 539 448
rect 533 445 539 446
rect 552 448 558 449
rect 552 446 554 448
rect 556 446 558 448
rect 552 445 558 446
rect 604 445 610 451
rect 17 428 23 429
rect 17 426 19 428
rect 21 426 23 428
rect 17 425 23 426
rect 36 428 42 429
rect 36 426 38 428
rect 40 426 42 428
rect 36 425 42 426
rect 109 423 115 429
rect 71 422 91 423
rect 71 420 87 422
rect 89 420 91 422
rect 109 421 111 423
rect 113 421 115 423
rect 109 420 115 421
rect 122 420 126 422
rect 71 419 91 420
rect 14 415 32 416
rect 14 413 28 415
rect 30 413 32 415
rect 14 412 32 413
rect 14 406 18 412
rect 14 404 15 406
rect 17 404 18 406
rect 10 383 11 394
rect 14 391 18 404
rect 33 399 39 400
rect 59 416 60 418
rect 71 415 75 419
rect 122 418 123 420
rect 125 418 126 420
rect 63 411 75 415
rect 63 406 67 411
rect 63 404 64 406
rect 66 404 67 406
rect 14 387 29 391
rect 25 383 29 387
rect 63 392 67 404
rect 96 415 100 417
rect 96 413 97 415
rect 99 413 100 415
rect 96 407 100 413
rect 122 415 126 418
rect 122 411 146 415
rect 96 403 107 407
rect 63 389 80 392
rect 63 388 77 389
rect 76 387 77 388
rect 79 387 80 389
rect 65 384 71 385
rect 25 382 42 383
rect 25 380 38 382
rect 40 380 42 382
rect 25 379 42 380
rect 65 382 67 384
rect 69 382 71 384
rect 17 375 23 376
rect 17 373 19 375
rect 21 373 23 375
rect 65 373 71 382
rect 76 382 80 387
rect 103 397 107 403
rect 142 407 146 411
rect 122 406 138 407
rect 122 404 134 406
rect 136 404 138 406
rect 122 403 138 404
rect 142 405 147 407
rect 142 403 144 405
rect 146 403 147 405
rect 122 397 126 403
rect 142 401 147 403
rect 142 399 146 401
rect 103 396 126 397
rect 103 394 105 396
rect 107 394 126 396
rect 103 393 126 394
rect 76 380 77 382
rect 79 380 80 382
rect 76 378 80 380
rect 85 382 91 383
rect 85 380 87 382
rect 89 380 91 382
rect 85 373 91 380
rect 114 382 118 384
rect 114 380 115 382
rect 117 380 118 382
rect 114 375 118 380
rect 122 382 126 393
rect 130 396 146 399
rect 130 394 131 396
rect 133 395 146 396
rect 133 394 134 395
rect 130 389 134 394
rect 130 387 131 389
rect 133 387 134 389
rect 130 385 134 387
rect 223 423 229 429
rect 185 422 205 423
rect 185 420 201 422
rect 203 420 205 422
rect 223 421 225 423
rect 227 421 229 423
rect 223 420 229 421
rect 236 420 240 422
rect 185 419 205 420
rect 173 416 174 418
rect 185 415 189 419
rect 236 418 237 420
rect 239 418 240 420
rect 280 422 300 423
rect 280 420 282 422
rect 284 420 300 422
rect 280 419 300 420
rect 177 411 189 415
rect 177 406 181 411
rect 177 404 178 406
rect 180 404 181 406
rect 177 392 181 404
rect 210 415 214 417
rect 210 413 211 415
rect 213 413 214 415
rect 210 407 214 413
rect 236 415 240 418
rect 236 411 260 415
rect 210 403 221 407
rect 177 389 194 392
rect 177 388 191 389
rect 190 387 191 388
rect 193 387 194 389
rect 179 384 185 385
rect 179 382 181 384
rect 183 382 185 384
rect 122 381 155 382
rect 122 379 151 381
rect 153 379 155 381
rect 122 378 155 379
rect 114 373 115 375
rect 117 373 118 375
rect 179 373 185 382
rect 190 382 194 387
rect 217 397 221 403
rect 256 407 260 411
rect 236 406 252 407
rect 236 404 248 406
rect 250 404 252 406
rect 236 403 252 404
rect 256 405 261 407
rect 256 403 258 405
rect 260 403 261 405
rect 236 397 240 403
rect 256 401 261 403
rect 256 399 260 401
rect 217 396 240 397
rect 217 394 219 396
rect 221 394 240 396
rect 217 393 240 394
rect 190 380 191 382
rect 193 380 194 382
rect 190 378 194 380
rect 199 382 205 383
rect 199 380 201 382
rect 203 380 205 382
rect 199 373 205 380
rect 228 382 232 384
rect 228 380 229 382
rect 231 380 232 382
rect 228 375 232 380
rect 236 382 240 393
rect 244 396 260 399
rect 244 394 245 396
rect 247 395 260 396
rect 296 415 300 419
rect 311 416 312 418
rect 296 411 308 415
rect 304 406 308 411
rect 304 404 305 406
rect 307 404 308 406
rect 247 394 248 395
rect 244 389 248 394
rect 244 387 245 389
rect 247 387 248 389
rect 244 385 248 387
rect 304 392 308 404
rect 291 389 308 392
rect 291 387 292 389
rect 294 388 308 389
rect 322 421 328 422
rect 322 419 324 421
rect 326 419 328 421
rect 322 418 328 419
rect 332 421 338 429
rect 332 419 334 421
rect 336 419 338 421
rect 349 423 364 424
rect 349 421 351 423
rect 353 421 364 423
rect 349 420 364 421
rect 332 418 338 419
rect 322 398 326 418
rect 360 415 364 420
rect 367 423 371 429
rect 367 421 368 423
rect 370 421 371 423
rect 367 419 371 421
rect 346 412 357 414
rect 346 410 354 412
rect 356 410 357 412
rect 360 413 374 415
rect 360 411 375 413
rect 346 408 357 410
rect 370 409 372 411
rect 374 409 375 411
rect 346 398 350 408
rect 370 407 375 409
rect 322 397 350 398
rect 322 395 324 397
rect 326 396 350 397
rect 326 395 347 396
rect 322 394 347 395
rect 349 394 350 396
rect 366 397 367 403
rect 346 392 350 394
rect 294 387 295 388
rect 280 382 286 383
rect 236 381 269 382
rect 236 379 265 381
rect 267 379 269 381
rect 236 378 269 379
rect 280 380 282 382
rect 284 380 286 382
rect 228 373 229 375
rect 231 373 232 375
rect 280 373 286 380
rect 291 382 295 387
rect 370 390 374 407
rect 358 386 374 390
rect 291 380 292 382
rect 294 380 295 382
rect 291 378 295 380
rect 300 384 306 385
rect 300 382 302 384
rect 304 382 306 384
rect 300 373 306 382
rect 349 385 362 386
rect 349 383 351 385
rect 353 383 362 385
rect 349 382 362 383
rect 400 423 404 429
rect 400 421 401 423
rect 403 421 404 423
rect 400 419 404 421
rect 407 423 422 424
rect 407 421 418 423
rect 420 421 422 423
rect 407 420 422 421
rect 433 421 439 429
rect 467 423 471 429
rect 407 415 411 420
rect 433 419 435 421
rect 437 419 439 421
rect 433 418 439 419
rect 443 421 449 422
rect 443 419 445 421
rect 447 419 449 421
rect 443 418 449 419
rect 397 413 411 415
rect 396 411 411 413
rect 414 412 425 414
rect 396 409 397 411
rect 399 409 401 411
rect 396 407 401 409
rect 414 410 415 412
rect 417 410 425 412
rect 414 408 425 410
rect 397 390 401 407
rect 404 397 405 403
rect 421 398 425 408
rect 445 398 449 418
rect 421 397 449 398
rect 421 396 445 397
rect 421 394 422 396
rect 424 395 445 396
rect 447 395 449 397
rect 424 394 449 395
rect 467 421 468 423
rect 470 421 471 423
rect 467 419 471 421
rect 474 423 489 424
rect 474 421 485 423
rect 487 421 489 423
rect 474 420 489 421
rect 500 421 506 429
rect 533 428 539 429
rect 533 426 535 428
rect 537 426 539 428
rect 533 425 539 426
rect 552 428 558 429
rect 552 426 554 428
rect 556 426 558 428
rect 552 425 558 426
rect 604 423 610 429
rect 474 415 478 420
rect 500 419 502 421
rect 504 419 506 421
rect 500 418 506 419
rect 510 421 516 422
rect 510 419 512 421
rect 514 419 516 421
rect 510 418 516 419
rect 464 413 478 415
rect 421 392 425 394
rect 397 386 413 390
rect 409 385 422 386
rect 409 383 418 385
rect 420 383 422 385
rect 409 382 422 383
rect 463 411 478 413
rect 481 412 492 414
rect 463 409 464 411
rect 466 409 468 411
rect 463 407 468 409
rect 481 410 482 412
rect 484 410 492 412
rect 481 408 492 410
rect 464 390 468 407
rect 471 397 472 403
rect 488 398 492 408
rect 512 398 516 418
rect 593 420 597 422
rect 604 421 606 423
rect 608 421 610 423
rect 604 420 610 421
rect 488 397 516 398
rect 488 396 512 397
rect 488 394 489 396
rect 491 395 512 396
rect 514 395 516 397
rect 491 394 516 395
rect 530 415 548 416
rect 530 413 544 415
rect 546 413 548 415
rect 530 412 548 413
rect 488 392 492 394
rect 530 406 534 412
rect 530 404 531 406
rect 533 404 534 406
rect 464 386 480 390
rect 476 385 489 386
rect 476 383 485 385
rect 487 383 489 385
rect 476 382 489 383
rect 526 383 527 394
rect 530 391 534 404
rect 593 418 594 420
rect 596 418 597 420
rect 593 415 597 418
rect 549 399 555 400
rect 530 387 545 391
rect 541 383 545 387
rect 573 411 597 415
rect 573 407 577 411
rect 619 415 623 417
rect 619 413 620 415
rect 622 413 623 415
rect 572 405 577 407
rect 572 403 573 405
rect 575 403 577 405
rect 581 406 597 407
rect 581 404 583 406
rect 585 404 597 406
rect 581 403 597 404
rect 572 401 577 403
rect 573 399 577 401
rect 573 396 589 399
rect 573 395 586 396
rect 585 394 586 395
rect 588 394 589 396
rect 585 389 589 394
rect 585 387 586 389
rect 588 387 589 389
rect 585 385 589 387
rect 593 397 597 403
rect 619 407 623 413
rect 612 403 623 407
rect 612 397 616 403
rect 593 396 616 397
rect 593 394 612 396
rect 614 394 616 396
rect 593 393 616 394
rect 541 382 558 383
rect 593 382 597 393
rect 541 380 554 382
rect 556 380 558 382
rect 541 379 558 380
rect 564 381 597 382
rect 564 379 566 381
rect 568 379 597 381
rect 564 378 597 379
rect 601 382 605 384
rect 601 380 602 382
rect 604 380 605 382
rect 333 375 337 377
rect 333 373 334 375
rect 336 373 337 375
rect 366 375 372 376
rect 366 373 368 375
rect 370 373 372 375
rect 399 375 405 376
rect 399 373 401 375
rect 403 373 405 375
rect 434 375 438 377
rect 434 373 435 375
rect 437 373 438 375
rect 466 375 472 376
rect 466 373 468 375
rect 470 373 472 375
rect 501 375 505 377
rect 501 373 502 375
rect 504 373 505 375
rect 533 375 539 376
rect 533 373 535 375
rect 537 373 539 375
rect 601 375 605 380
rect 601 373 602 375
rect 604 373 605 375
rect 17 355 19 357
rect 21 355 23 357
rect 17 354 23 355
rect 25 350 42 351
rect 25 348 38 350
rect 40 348 42 350
rect 25 347 42 348
rect 65 348 71 357
rect 10 336 11 347
rect 25 343 29 347
rect 65 346 67 348
rect 69 346 71 348
rect 65 345 71 346
rect 76 350 80 352
rect 76 348 77 350
rect 79 348 80 350
rect 14 339 29 343
rect 76 343 80 348
rect 85 350 91 357
rect 114 355 115 357
rect 117 355 118 357
rect 85 348 87 350
rect 89 348 91 350
rect 85 347 91 348
rect 114 350 118 355
rect 114 348 115 350
rect 117 348 118 350
rect 114 346 118 348
rect 122 351 155 352
rect 122 349 151 351
rect 153 349 155 351
rect 122 348 155 349
rect 179 348 185 357
rect 76 342 77 343
rect 14 326 18 339
rect 63 341 77 342
rect 79 341 80 343
rect 63 338 80 341
rect 33 330 39 331
rect 14 324 15 326
rect 17 324 18 326
rect 14 318 18 324
rect 14 317 32 318
rect 14 315 28 317
rect 30 315 32 317
rect 14 314 32 315
rect 63 326 67 338
rect 122 337 126 348
rect 179 346 181 348
rect 183 346 185 348
rect 179 345 185 346
rect 190 350 194 352
rect 190 348 191 350
rect 193 348 194 350
rect 103 336 126 337
rect 103 334 105 336
rect 107 334 126 336
rect 103 333 126 334
rect 103 327 107 333
rect 63 324 64 326
rect 66 324 67 326
rect 63 319 67 324
rect 63 315 75 319
rect 59 312 60 314
rect 71 311 75 315
rect 96 323 107 327
rect 96 317 100 323
rect 122 327 126 333
rect 130 343 134 345
rect 130 341 131 343
rect 133 341 134 343
rect 130 336 134 341
rect 130 334 131 336
rect 133 335 134 336
rect 133 334 146 335
rect 130 331 146 334
rect 142 329 146 331
rect 142 327 147 329
rect 122 326 138 327
rect 122 324 134 326
rect 136 324 138 326
rect 122 323 138 324
rect 142 325 144 327
rect 146 325 147 327
rect 142 323 147 325
rect 96 315 97 317
rect 99 315 100 317
rect 96 313 100 315
rect 142 319 146 323
rect 122 315 146 319
rect 122 312 126 315
rect 71 310 91 311
rect 122 310 123 312
rect 125 310 126 312
rect 71 308 87 310
rect 89 308 91 310
rect 71 307 91 308
rect 109 309 115 310
rect 109 307 111 309
rect 113 307 115 309
rect 122 308 126 310
rect 190 343 194 348
rect 199 350 205 357
rect 228 355 229 357
rect 231 355 232 357
rect 199 348 201 350
rect 203 348 205 350
rect 199 347 205 348
rect 228 350 232 355
rect 228 348 229 350
rect 231 348 232 350
rect 228 346 232 348
rect 236 351 269 352
rect 236 349 265 351
rect 267 349 269 351
rect 236 348 269 349
rect 280 350 286 357
rect 280 348 282 350
rect 284 348 286 350
rect 190 342 191 343
rect 177 341 191 342
rect 193 341 194 343
rect 177 338 194 341
rect 177 326 181 338
rect 236 337 240 348
rect 280 347 286 348
rect 291 350 295 352
rect 291 348 292 350
rect 294 348 295 350
rect 217 336 240 337
rect 217 334 219 336
rect 221 334 240 336
rect 217 333 240 334
rect 217 327 221 333
rect 177 324 178 326
rect 180 324 181 326
rect 177 319 181 324
rect 177 315 189 319
rect 173 312 174 314
rect 17 304 23 305
rect 17 302 19 304
rect 21 302 23 304
rect 17 301 23 302
rect 36 304 42 305
rect 36 302 38 304
rect 40 302 42 304
rect 36 301 42 302
rect 109 301 115 307
rect 185 311 189 315
rect 210 323 221 327
rect 210 317 214 323
rect 236 327 240 333
rect 244 343 248 345
rect 244 341 245 343
rect 247 341 248 343
rect 244 336 248 341
rect 244 334 245 336
rect 247 335 248 336
rect 247 334 260 335
rect 244 331 260 334
rect 256 329 260 331
rect 291 343 295 348
rect 300 348 306 357
rect 333 355 334 357
rect 336 355 337 357
rect 333 353 337 355
rect 366 355 368 357
rect 370 355 372 357
rect 366 354 372 355
rect 399 355 401 357
rect 403 355 405 357
rect 399 354 405 355
rect 434 355 435 357
rect 437 355 438 357
rect 434 353 438 355
rect 466 355 468 357
rect 470 355 472 357
rect 466 354 472 355
rect 501 355 502 357
rect 504 355 505 357
rect 501 353 505 355
rect 533 355 535 357
rect 537 355 539 357
rect 533 354 539 355
rect 601 355 602 357
rect 604 355 605 357
rect 300 346 302 348
rect 304 346 306 348
rect 300 345 306 346
rect 291 341 292 343
rect 294 342 295 343
rect 294 341 308 342
rect 291 338 308 341
rect 256 327 261 329
rect 236 326 252 327
rect 236 324 248 326
rect 250 324 252 326
rect 236 323 252 324
rect 256 325 258 327
rect 260 325 261 327
rect 256 323 261 325
rect 210 315 211 317
rect 213 315 214 317
rect 210 313 214 315
rect 256 319 260 323
rect 236 315 260 319
rect 236 312 240 315
rect 185 310 205 311
rect 236 310 237 312
rect 239 310 240 312
rect 304 326 308 338
rect 349 347 362 348
rect 349 345 351 347
rect 353 345 362 347
rect 349 344 362 345
rect 358 340 374 344
rect 346 336 350 338
rect 304 324 305 326
rect 307 324 308 326
rect 304 319 308 324
rect 296 315 308 319
rect 296 311 300 315
rect 311 312 312 314
rect 185 308 201 310
rect 203 308 205 310
rect 185 307 205 308
rect 223 309 229 310
rect 223 307 225 309
rect 227 307 229 309
rect 236 308 240 310
rect 280 310 300 311
rect 280 308 282 310
rect 284 308 300 310
rect 280 307 300 308
rect 223 301 229 307
rect 322 335 347 336
rect 322 333 324 335
rect 326 334 347 335
rect 349 334 350 336
rect 326 333 350 334
rect 322 332 350 333
rect 322 312 326 332
rect 346 322 350 332
rect 366 327 367 333
rect 370 323 374 340
rect 346 320 357 322
rect 346 318 354 320
rect 356 318 357 320
rect 370 321 375 323
rect 370 319 372 321
rect 374 319 375 321
rect 346 316 357 318
rect 360 317 375 319
rect 360 315 374 317
rect 322 311 328 312
rect 322 309 324 311
rect 326 309 328 311
rect 322 308 328 309
rect 332 311 338 312
rect 332 309 334 311
rect 336 309 338 311
rect 360 310 364 315
rect 332 301 338 309
rect 349 309 364 310
rect 349 307 351 309
rect 353 307 364 309
rect 349 306 364 307
rect 367 309 371 311
rect 367 307 368 309
rect 370 307 371 309
rect 367 301 371 307
rect 409 347 422 348
rect 409 345 418 347
rect 420 345 422 347
rect 409 344 422 345
rect 397 340 413 344
rect 397 323 401 340
rect 476 347 489 348
rect 421 336 425 338
rect 404 327 405 333
rect 421 334 422 336
rect 424 335 449 336
rect 424 334 445 335
rect 421 333 445 334
rect 447 333 449 335
rect 421 332 449 333
rect 396 321 401 323
rect 421 322 425 332
rect 396 319 397 321
rect 399 319 401 321
rect 414 320 425 322
rect 396 317 411 319
rect 397 315 411 317
rect 414 318 415 320
rect 417 318 425 320
rect 414 316 425 318
rect 400 309 404 311
rect 400 307 401 309
rect 403 307 404 309
rect 400 301 404 307
rect 407 310 411 315
rect 445 312 449 332
rect 433 311 439 312
rect 407 309 422 310
rect 407 307 418 309
rect 420 307 422 309
rect 407 306 422 307
rect 433 309 435 311
rect 437 309 439 311
rect 433 301 439 309
rect 443 311 449 312
rect 443 309 445 311
rect 447 309 449 311
rect 443 308 449 309
rect 476 345 485 347
rect 487 345 489 347
rect 476 344 489 345
rect 464 340 480 344
rect 464 323 468 340
rect 564 351 597 352
rect 541 350 558 351
rect 541 348 554 350
rect 556 348 558 350
rect 564 349 566 351
rect 568 349 597 351
rect 564 348 597 349
rect 541 347 558 348
rect 488 336 492 338
rect 471 327 472 333
rect 488 334 489 336
rect 491 335 516 336
rect 491 334 512 335
rect 488 333 512 334
rect 514 333 516 335
rect 488 332 516 333
rect 463 321 468 323
rect 488 322 492 332
rect 463 319 464 321
rect 466 319 468 321
rect 481 320 492 322
rect 463 317 478 319
rect 464 315 478 317
rect 481 318 482 320
rect 484 318 492 320
rect 481 316 492 318
rect 467 309 471 311
rect 467 307 468 309
rect 470 307 471 309
rect 467 301 471 307
rect 474 310 478 315
rect 512 312 516 332
rect 526 336 527 347
rect 541 343 545 347
rect 530 339 545 343
rect 530 326 534 339
rect 585 343 589 345
rect 585 341 586 343
rect 588 341 589 343
rect 549 330 555 331
rect 530 324 531 326
rect 533 324 534 326
rect 530 318 534 324
rect 530 317 548 318
rect 530 315 544 317
rect 546 315 548 317
rect 530 314 548 315
rect 585 336 589 341
rect 585 335 586 336
rect 573 334 586 335
rect 588 334 589 336
rect 573 331 589 334
rect 593 337 597 348
rect 601 350 605 355
rect 601 348 602 350
rect 604 348 605 350
rect 601 346 605 348
rect 593 336 616 337
rect 593 334 612 336
rect 614 334 616 336
rect 593 333 616 334
rect 573 329 577 331
rect 572 327 577 329
rect 593 327 597 333
rect 572 325 573 327
rect 575 325 577 327
rect 572 323 577 325
rect 581 326 597 327
rect 581 324 583 326
rect 585 324 597 326
rect 581 323 597 324
rect 500 311 506 312
rect 474 309 489 310
rect 474 307 485 309
rect 487 307 489 309
rect 474 306 489 307
rect 500 309 502 311
rect 504 309 506 311
rect 500 301 506 309
rect 510 311 516 312
rect 510 309 512 311
rect 514 309 516 311
rect 510 308 516 309
rect 573 319 577 323
rect 612 327 616 333
rect 612 323 623 327
rect 573 315 597 319
rect 593 312 597 315
rect 619 317 623 323
rect 619 315 620 317
rect 622 315 623 317
rect 619 313 623 315
rect 593 310 594 312
rect 596 310 597 312
rect 593 308 597 310
rect 604 309 610 310
rect 604 307 606 309
rect 608 307 610 309
rect 533 304 539 305
rect 533 302 535 304
rect 537 302 539 304
rect 533 301 539 302
rect 552 304 558 305
rect 552 302 554 304
rect 556 302 558 304
rect 552 301 558 302
rect 604 301 610 307
rect 17 284 23 285
rect 17 282 19 284
rect 21 282 23 284
rect 17 281 23 282
rect 36 284 42 285
rect 36 282 38 284
rect 40 282 42 284
rect 36 281 42 282
rect 109 279 115 285
rect 71 278 91 279
rect 71 276 87 278
rect 89 276 91 278
rect 109 277 111 279
rect 113 277 115 279
rect 109 276 115 277
rect 122 276 126 278
rect 71 275 91 276
rect 14 271 32 272
rect 14 269 28 271
rect 30 269 32 271
rect 14 268 32 269
rect 14 262 18 268
rect 14 260 15 262
rect 17 260 18 262
rect 10 239 11 250
rect 14 247 18 260
rect 33 255 39 256
rect 59 272 60 274
rect 71 271 75 275
rect 122 274 123 276
rect 125 274 126 276
rect 63 267 75 271
rect 63 262 67 267
rect 63 260 64 262
rect 66 260 67 262
rect 14 243 29 247
rect 25 239 29 243
rect 63 248 67 260
rect 96 271 100 273
rect 96 269 97 271
rect 99 269 100 271
rect 96 263 100 269
rect 122 271 126 274
rect 122 267 146 271
rect 96 259 107 263
rect 63 245 80 248
rect 63 244 77 245
rect 76 243 77 244
rect 79 243 80 245
rect 65 240 71 241
rect 25 238 42 239
rect 25 236 38 238
rect 40 236 42 238
rect 25 235 42 236
rect 65 238 67 240
rect 69 238 71 240
rect 17 231 23 232
rect 17 229 19 231
rect 21 229 23 231
rect 65 229 71 238
rect 76 238 80 243
rect 103 253 107 259
rect 142 263 146 267
rect 122 262 138 263
rect 122 260 134 262
rect 136 260 138 262
rect 122 259 138 260
rect 142 261 147 263
rect 142 259 144 261
rect 146 259 147 261
rect 122 253 126 259
rect 142 257 147 259
rect 142 255 146 257
rect 103 252 126 253
rect 103 250 105 252
rect 107 250 126 252
rect 103 249 126 250
rect 76 236 77 238
rect 79 236 80 238
rect 76 234 80 236
rect 85 238 91 239
rect 85 236 87 238
rect 89 236 91 238
rect 85 229 91 236
rect 114 238 118 240
rect 114 236 115 238
rect 117 236 118 238
rect 114 231 118 236
rect 122 238 126 249
rect 130 252 146 255
rect 130 250 131 252
rect 133 251 146 252
rect 133 250 134 251
rect 130 245 134 250
rect 130 243 131 245
rect 133 243 134 245
rect 130 241 134 243
rect 223 279 229 285
rect 185 278 205 279
rect 185 276 201 278
rect 203 276 205 278
rect 223 277 225 279
rect 227 277 229 279
rect 223 276 229 277
rect 236 276 240 278
rect 185 275 205 276
rect 173 272 174 274
rect 185 271 189 275
rect 236 274 237 276
rect 239 274 240 276
rect 280 278 300 279
rect 280 276 282 278
rect 284 276 300 278
rect 280 275 300 276
rect 177 267 189 271
rect 177 262 181 267
rect 177 260 178 262
rect 180 260 181 262
rect 177 248 181 260
rect 210 271 214 273
rect 210 269 211 271
rect 213 269 214 271
rect 210 263 214 269
rect 236 271 240 274
rect 236 267 260 271
rect 210 259 221 263
rect 177 245 194 248
rect 177 244 191 245
rect 190 243 191 244
rect 193 243 194 245
rect 179 240 185 241
rect 179 238 181 240
rect 183 238 185 240
rect 122 237 155 238
rect 122 235 151 237
rect 153 235 155 237
rect 122 234 155 235
rect 114 229 115 231
rect 117 229 118 231
rect 179 229 185 238
rect 190 238 194 243
rect 217 253 221 259
rect 256 263 260 267
rect 236 262 252 263
rect 236 260 248 262
rect 250 260 252 262
rect 236 259 252 260
rect 256 261 261 263
rect 256 259 258 261
rect 260 259 261 261
rect 236 253 240 259
rect 256 257 261 259
rect 256 255 260 257
rect 217 252 240 253
rect 217 250 219 252
rect 221 250 240 252
rect 217 249 240 250
rect 190 236 191 238
rect 193 236 194 238
rect 190 234 194 236
rect 199 238 205 239
rect 199 236 201 238
rect 203 236 205 238
rect 199 229 205 236
rect 228 238 232 240
rect 228 236 229 238
rect 231 236 232 238
rect 228 231 232 236
rect 236 238 240 249
rect 244 252 260 255
rect 244 250 245 252
rect 247 251 260 252
rect 296 271 300 275
rect 311 272 312 274
rect 296 267 308 271
rect 304 262 308 267
rect 304 260 305 262
rect 307 260 308 262
rect 247 250 248 251
rect 244 245 248 250
rect 244 243 245 245
rect 247 243 248 245
rect 244 241 248 243
rect 304 248 308 260
rect 291 245 308 248
rect 291 243 292 245
rect 294 244 308 245
rect 322 277 328 278
rect 322 275 324 277
rect 326 275 328 277
rect 322 274 328 275
rect 332 277 338 285
rect 332 275 334 277
rect 336 275 338 277
rect 349 279 364 280
rect 349 277 351 279
rect 353 277 364 279
rect 349 276 364 277
rect 332 274 338 275
rect 322 254 326 274
rect 360 271 364 276
rect 367 279 371 285
rect 367 277 368 279
rect 370 277 371 279
rect 367 275 371 277
rect 346 268 357 270
rect 346 266 354 268
rect 356 266 357 268
rect 360 269 374 271
rect 360 267 375 269
rect 346 264 357 266
rect 370 265 372 267
rect 374 265 375 267
rect 346 254 350 264
rect 370 263 375 265
rect 322 253 350 254
rect 322 251 324 253
rect 326 252 350 253
rect 326 251 347 252
rect 322 250 347 251
rect 349 250 350 252
rect 366 253 367 259
rect 346 248 350 250
rect 294 243 295 244
rect 280 238 286 239
rect 236 237 269 238
rect 236 235 265 237
rect 267 235 269 237
rect 236 234 269 235
rect 280 236 282 238
rect 284 236 286 238
rect 228 229 229 231
rect 231 229 232 231
rect 280 229 286 236
rect 291 238 295 243
rect 370 246 374 263
rect 358 242 374 246
rect 291 236 292 238
rect 294 236 295 238
rect 291 234 295 236
rect 300 240 306 241
rect 300 238 302 240
rect 304 238 306 240
rect 300 229 306 238
rect 349 241 362 242
rect 349 239 351 241
rect 353 239 362 241
rect 349 238 362 239
rect 400 279 404 285
rect 400 277 401 279
rect 403 277 404 279
rect 400 275 404 277
rect 407 279 422 280
rect 407 277 418 279
rect 420 277 422 279
rect 407 276 422 277
rect 433 277 439 285
rect 467 279 471 285
rect 407 271 411 276
rect 433 275 435 277
rect 437 275 439 277
rect 433 274 439 275
rect 443 277 449 278
rect 443 275 445 277
rect 447 275 449 277
rect 443 274 449 275
rect 397 269 411 271
rect 396 267 411 269
rect 414 268 425 270
rect 396 265 397 267
rect 399 265 401 267
rect 396 263 401 265
rect 414 266 415 268
rect 417 266 425 268
rect 414 264 425 266
rect 397 246 401 263
rect 404 253 405 259
rect 421 254 425 264
rect 445 254 449 274
rect 421 253 449 254
rect 421 252 445 253
rect 421 250 422 252
rect 424 251 445 252
rect 447 251 449 253
rect 424 250 449 251
rect 467 277 468 279
rect 470 277 471 279
rect 467 275 471 277
rect 474 279 489 280
rect 474 277 485 279
rect 487 277 489 279
rect 474 276 489 277
rect 500 277 506 285
rect 533 284 539 285
rect 533 282 535 284
rect 537 282 539 284
rect 533 281 539 282
rect 552 284 558 285
rect 552 282 554 284
rect 556 282 558 284
rect 552 281 558 282
rect 604 279 610 285
rect 474 271 478 276
rect 500 275 502 277
rect 504 275 506 277
rect 500 274 506 275
rect 510 277 516 278
rect 510 275 512 277
rect 514 275 516 277
rect 510 274 516 275
rect 464 269 478 271
rect 421 248 425 250
rect 397 242 413 246
rect 409 241 422 242
rect 409 239 418 241
rect 420 239 422 241
rect 409 238 422 239
rect 463 267 478 269
rect 481 268 492 270
rect 463 265 464 267
rect 466 265 468 267
rect 463 263 468 265
rect 481 266 482 268
rect 484 266 492 268
rect 481 264 492 266
rect 464 246 468 263
rect 471 253 472 259
rect 488 254 492 264
rect 512 254 516 274
rect 593 276 597 278
rect 604 277 606 279
rect 608 277 610 279
rect 604 276 610 277
rect 488 253 516 254
rect 488 252 512 253
rect 488 250 489 252
rect 491 251 512 252
rect 514 251 516 253
rect 491 250 516 251
rect 530 271 548 272
rect 530 269 544 271
rect 546 269 548 271
rect 530 268 548 269
rect 488 248 492 250
rect 530 262 534 268
rect 530 260 531 262
rect 533 260 534 262
rect 464 242 480 246
rect 476 241 489 242
rect 476 239 485 241
rect 487 239 489 241
rect 476 238 489 239
rect 526 239 527 250
rect 530 247 534 260
rect 593 274 594 276
rect 596 274 597 276
rect 593 271 597 274
rect 549 255 555 256
rect 530 243 545 247
rect 541 239 545 243
rect 573 267 597 271
rect 573 263 577 267
rect 619 271 623 273
rect 619 269 620 271
rect 622 269 623 271
rect 572 261 577 263
rect 572 259 573 261
rect 575 259 577 261
rect 581 262 597 263
rect 581 260 583 262
rect 585 260 597 262
rect 581 259 597 260
rect 572 257 577 259
rect 573 255 577 257
rect 573 252 589 255
rect 573 251 586 252
rect 585 250 586 251
rect 588 250 589 252
rect 585 245 589 250
rect 585 243 586 245
rect 588 243 589 245
rect 585 241 589 243
rect 593 253 597 259
rect 619 263 623 269
rect 612 259 623 263
rect 612 253 616 259
rect 593 252 616 253
rect 593 250 612 252
rect 614 250 616 252
rect 593 249 616 250
rect 541 238 558 239
rect 593 238 597 249
rect 541 236 554 238
rect 556 236 558 238
rect 541 235 558 236
rect 564 237 597 238
rect 564 235 566 237
rect 568 235 597 237
rect 564 234 597 235
rect 601 238 605 240
rect 601 236 602 238
rect 604 236 605 238
rect 333 231 337 233
rect 333 229 334 231
rect 336 229 337 231
rect 366 231 372 232
rect 366 229 368 231
rect 370 229 372 231
rect 399 231 405 232
rect 399 229 401 231
rect 403 229 405 231
rect 434 231 438 233
rect 434 229 435 231
rect 437 229 438 231
rect 466 231 472 232
rect 466 229 468 231
rect 470 229 472 231
rect 501 231 505 233
rect 501 229 502 231
rect 504 229 505 231
rect 533 231 539 232
rect 533 229 535 231
rect 537 229 539 231
rect 601 231 605 236
rect 601 229 602 231
rect 604 229 605 231
rect 17 211 19 213
rect 21 211 23 213
rect 17 210 23 211
rect 25 206 42 207
rect 25 204 38 206
rect 40 204 42 206
rect 25 203 42 204
rect 65 204 71 213
rect 10 192 11 203
rect 25 199 29 203
rect 65 202 67 204
rect 69 202 71 204
rect 65 201 71 202
rect 76 206 80 208
rect 76 204 77 206
rect 79 204 80 206
rect 14 195 29 199
rect 76 199 80 204
rect 85 206 91 213
rect 114 211 115 213
rect 117 211 118 213
rect 85 204 87 206
rect 89 204 91 206
rect 85 203 91 204
rect 114 206 118 211
rect 114 204 115 206
rect 117 204 118 206
rect 114 202 118 204
rect 122 207 155 208
rect 122 205 151 207
rect 153 205 155 207
rect 122 204 155 205
rect 179 204 185 213
rect 76 198 77 199
rect 14 182 18 195
rect 63 197 77 198
rect 79 197 80 199
rect 63 194 80 197
rect 33 186 39 187
rect 14 180 15 182
rect 17 180 18 182
rect 14 174 18 180
rect 14 173 32 174
rect 14 171 28 173
rect 30 171 32 173
rect 14 170 32 171
rect 63 182 67 194
rect 122 193 126 204
rect 179 202 181 204
rect 183 202 185 204
rect 179 201 185 202
rect 190 206 194 208
rect 190 204 191 206
rect 193 204 194 206
rect 103 192 126 193
rect 103 190 105 192
rect 107 190 126 192
rect 103 189 126 190
rect 103 183 107 189
rect 63 180 64 182
rect 66 180 67 182
rect 63 175 67 180
rect 63 171 75 175
rect 59 168 60 170
rect 71 167 75 171
rect 96 179 107 183
rect 96 173 100 179
rect 122 183 126 189
rect 130 199 134 201
rect 130 197 131 199
rect 133 197 134 199
rect 130 192 134 197
rect 130 190 131 192
rect 133 191 134 192
rect 133 190 146 191
rect 130 187 146 190
rect 142 185 146 187
rect 142 183 147 185
rect 122 182 138 183
rect 122 180 134 182
rect 136 180 138 182
rect 122 179 138 180
rect 142 181 144 183
rect 146 181 147 183
rect 142 179 147 181
rect 96 171 97 173
rect 99 171 100 173
rect 96 169 100 171
rect 142 175 146 179
rect 122 171 146 175
rect 122 168 126 171
rect 71 166 91 167
rect 122 166 123 168
rect 125 166 126 168
rect 71 164 87 166
rect 89 164 91 166
rect 71 163 91 164
rect 109 165 115 166
rect 109 163 111 165
rect 113 163 115 165
rect 122 164 126 166
rect 190 199 194 204
rect 199 206 205 213
rect 228 211 229 213
rect 231 211 232 213
rect 199 204 201 206
rect 203 204 205 206
rect 199 203 205 204
rect 228 206 232 211
rect 228 204 229 206
rect 231 204 232 206
rect 228 202 232 204
rect 236 207 269 208
rect 236 205 265 207
rect 267 205 269 207
rect 236 204 269 205
rect 280 206 286 213
rect 280 204 282 206
rect 284 204 286 206
rect 190 198 191 199
rect 177 197 191 198
rect 193 197 194 199
rect 177 194 194 197
rect 177 182 181 194
rect 236 193 240 204
rect 280 203 286 204
rect 291 206 295 208
rect 291 204 292 206
rect 294 204 295 206
rect 217 192 240 193
rect 217 190 219 192
rect 221 190 240 192
rect 217 189 240 190
rect 217 183 221 189
rect 177 180 178 182
rect 180 180 181 182
rect 177 175 181 180
rect 177 171 189 175
rect 173 168 174 170
rect 17 160 23 161
rect 17 158 19 160
rect 21 158 23 160
rect 17 157 23 158
rect 36 160 42 161
rect 36 158 38 160
rect 40 158 42 160
rect 36 157 42 158
rect 109 157 115 163
rect 185 167 189 171
rect 210 179 221 183
rect 210 173 214 179
rect 236 183 240 189
rect 244 199 248 201
rect 244 197 245 199
rect 247 197 248 199
rect 244 192 248 197
rect 244 190 245 192
rect 247 191 248 192
rect 247 190 260 191
rect 244 187 260 190
rect 256 185 260 187
rect 291 199 295 204
rect 300 204 306 213
rect 333 211 334 213
rect 336 211 337 213
rect 333 209 337 211
rect 366 211 368 213
rect 370 211 372 213
rect 366 210 372 211
rect 399 211 401 213
rect 403 211 405 213
rect 399 210 405 211
rect 434 211 435 213
rect 437 211 438 213
rect 434 209 438 211
rect 466 211 468 213
rect 470 211 472 213
rect 466 210 472 211
rect 501 211 502 213
rect 504 211 505 213
rect 501 209 505 211
rect 533 211 535 213
rect 537 211 539 213
rect 533 210 539 211
rect 601 211 602 213
rect 604 211 605 213
rect 300 202 302 204
rect 304 202 306 204
rect 300 201 306 202
rect 291 197 292 199
rect 294 198 295 199
rect 294 197 308 198
rect 291 194 308 197
rect 256 183 261 185
rect 236 182 252 183
rect 236 180 248 182
rect 250 180 252 182
rect 236 179 252 180
rect 256 181 258 183
rect 260 181 261 183
rect 256 179 261 181
rect 210 171 211 173
rect 213 171 214 173
rect 210 169 214 171
rect 256 175 260 179
rect 236 171 260 175
rect 236 168 240 171
rect 185 166 205 167
rect 236 166 237 168
rect 239 166 240 168
rect 304 182 308 194
rect 349 203 362 204
rect 349 201 351 203
rect 353 201 362 203
rect 349 200 362 201
rect 358 196 374 200
rect 346 192 350 194
rect 304 180 305 182
rect 307 180 308 182
rect 304 175 308 180
rect 296 171 308 175
rect 296 167 300 171
rect 311 168 312 170
rect 185 164 201 166
rect 203 164 205 166
rect 185 163 205 164
rect 223 165 229 166
rect 223 163 225 165
rect 227 163 229 165
rect 236 164 240 166
rect 280 166 300 167
rect 280 164 282 166
rect 284 164 300 166
rect 280 163 300 164
rect 223 157 229 163
rect 322 191 347 192
rect 322 189 324 191
rect 326 190 347 191
rect 349 190 350 192
rect 326 189 350 190
rect 322 188 350 189
rect 322 168 326 188
rect 346 178 350 188
rect 366 183 367 189
rect 370 179 374 196
rect 346 176 357 178
rect 346 174 354 176
rect 356 174 357 176
rect 370 177 375 179
rect 370 175 372 177
rect 374 175 375 177
rect 346 172 357 174
rect 360 173 375 175
rect 360 171 374 173
rect 322 167 328 168
rect 322 165 324 167
rect 326 165 328 167
rect 322 164 328 165
rect 332 167 338 168
rect 332 165 334 167
rect 336 165 338 167
rect 360 166 364 171
rect 332 157 338 165
rect 349 165 364 166
rect 349 163 351 165
rect 353 163 364 165
rect 349 162 364 163
rect 367 165 371 167
rect 367 163 368 165
rect 370 163 371 165
rect 367 157 371 163
rect 409 203 422 204
rect 409 201 418 203
rect 420 201 422 203
rect 409 200 422 201
rect 397 196 413 200
rect 397 179 401 196
rect 476 203 489 204
rect 421 192 425 194
rect 404 183 405 189
rect 421 190 422 192
rect 424 191 449 192
rect 424 190 445 191
rect 421 189 445 190
rect 447 189 449 191
rect 421 188 449 189
rect 396 177 401 179
rect 421 178 425 188
rect 396 175 397 177
rect 399 175 401 177
rect 414 176 425 178
rect 396 173 411 175
rect 397 171 411 173
rect 414 174 415 176
rect 417 174 425 176
rect 414 172 425 174
rect 400 165 404 167
rect 400 163 401 165
rect 403 163 404 165
rect 400 157 404 163
rect 407 166 411 171
rect 445 168 449 188
rect 433 167 439 168
rect 407 165 422 166
rect 407 163 418 165
rect 420 163 422 165
rect 407 162 422 163
rect 433 165 435 167
rect 437 165 439 167
rect 433 157 439 165
rect 443 167 449 168
rect 443 165 445 167
rect 447 165 449 167
rect 443 164 449 165
rect 476 201 485 203
rect 487 201 489 203
rect 476 200 489 201
rect 464 196 480 200
rect 464 179 468 196
rect 564 207 597 208
rect 541 206 558 207
rect 541 204 554 206
rect 556 204 558 206
rect 564 205 566 207
rect 568 205 597 207
rect 564 204 597 205
rect 541 203 558 204
rect 488 192 492 194
rect 471 183 472 189
rect 488 190 489 192
rect 491 191 516 192
rect 491 190 512 191
rect 488 189 512 190
rect 514 189 516 191
rect 488 188 516 189
rect 463 177 468 179
rect 488 178 492 188
rect 463 175 464 177
rect 466 175 468 177
rect 481 176 492 178
rect 463 173 478 175
rect 464 171 478 173
rect 481 174 482 176
rect 484 174 492 176
rect 481 172 492 174
rect 467 165 471 167
rect 467 163 468 165
rect 470 163 471 165
rect 467 157 471 163
rect 474 166 478 171
rect 512 168 516 188
rect 526 192 527 203
rect 541 199 545 203
rect 530 195 545 199
rect 530 182 534 195
rect 585 199 589 201
rect 585 197 586 199
rect 588 197 589 199
rect 549 186 555 187
rect 530 180 531 182
rect 533 180 534 182
rect 530 174 534 180
rect 530 173 548 174
rect 530 171 544 173
rect 546 171 548 173
rect 530 170 548 171
rect 585 192 589 197
rect 585 191 586 192
rect 573 190 586 191
rect 588 190 589 192
rect 573 187 589 190
rect 593 193 597 204
rect 601 206 605 211
rect 601 204 602 206
rect 604 204 605 206
rect 601 202 605 204
rect 593 192 616 193
rect 593 190 612 192
rect 614 190 616 192
rect 593 189 616 190
rect 573 185 577 187
rect 572 183 577 185
rect 593 183 597 189
rect 572 181 573 183
rect 575 181 577 183
rect 572 179 577 181
rect 581 182 597 183
rect 581 180 583 182
rect 585 180 597 182
rect 581 179 597 180
rect 500 167 506 168
rect 474 165 489 166
rect 474 163 485 165
rect 487 163 489 165
rect 474 162 489 163
rect 500 165 502 167
rect 504 165 506 167
rect 500 157 506 165
rect 510 167 516 168
rect 510 165 512 167
rect 514 165 516 167
rect 510 164 516 165
rect 573 175 577 179
rect 612 183 616 189
rect 612 179 623 183
rect 573 171 597 175
rect 593 168 597 171
rect 619 173 623 179
rect 619 171 620 173
rect 622 171 623 173
rect 619 169 623 171
rect 593 166 594 168
rect 596 166 597 168
rect 593 164 597 166
rect 604 165 610 166
rect 604 163 606 165
rect 608 163 610 165
rect 533 160 539 161
rect 533 158 535 160
rect 537 158 539 160
rect 533 157 539 158
rect 552 160 558 161
rect 552 158 554 160
rect 556 158 558 160
rect 552 157 558 158
rect 604 157 610 163
rect 17 140 23 141
rect 17 138 19 140
rect 21 138 23 140
rect 17 137 23 138
rect 36 140 42 141
rect 36 138 38 140
rect 40 138 42 140
rect 36 137 42 138
rect 109 135 115 141
rect 71 134 91 135
rect 71 132 87 134
rect 89 132 91 134
rect 109 133 111 135
rect 113 133 115 135
rect 109 132 115 133
rect 122 132 126 134
rect 71 131 91 132
rect 14 127 32 128
rect 14 125 28 127
rect 30 125 32 127
rect 14 124 32 125
rect 14 118 18 124
rect 14 116 15 118
rect 17 116 18 118
rect 10 95 11 106
rect 14 103 18 116
rect 33 111 39 112
rect 59 128 60 130
rect 71 127 75 131
rect 122 130 123 132
rect 125 130 126 132
rect 63 123 75 127
rect 63 118 67 123
rect 63 116 64 118
rect 66 116 67 118
rect 14 99 29 103
rect 25 95 29 99
rect 63 104 67 116
rect 96 127 100 129
rect 96 125 97 127
rect 99 125 100 127
rect 96 119 100 125
rect 122 127 126 130
rect 122 123 146 127
rect 96 115 107 119
rect 63 101 80 104
rect 63 100 77 101
rect 76 99 77 100
rect 79 99 80 101
rect 65 96 71 97
rect 25 94 42 95
rect 25 92 38 94
rect 40 92 42 94
rect 25 91 42 92
rect 65 94 67 96
rect 69 94 71 96
rect 17 87 23 88
rect 17 85 19 87
rect 21 85 23 87
rect 65 85 71 94
rect 76 94 80 99
rect 103 109 107 115
rect 142 119 146 123
rect 122 118 138 119
rect 122 116 134 118
rect 136 116 138 118
rect 122 115 138 116
rect 142 117 147 119
rect 142 115 144 117
rect 146 115 147 117
rect 122 109 126 115
rect 142 113 147 115
rect 142 111 146 113
rect 103 108 126 109
rect 103 106 105 108
rect 107 106 126 108
rect 103 105 126 106
rect 76 92 77 94
rect 79 92 80 94
rect 76 90 80 92
rect 85 94 91 95
rect 85 92 87 94
rect 89 92 91 94
rect 85 85 91 92
rect 114 94 118 96
rect 114 92 115 94
rect 117 92 118 94
rect 114 87 118 92
rect 122 94 126 105
rect 130 108 146 111
rect 130 106 131 108
rect 133 107 146 108
rect 133 106 134 107
rect 130 101 134 106
rect 130 99 131 101
rect 133 99 134 101
rect 130 97 134 99
rect 223 135 229 141
rect 185 134 205 135
rect 185 132 201 134
rect 203 132 205 134
rect 223 133 225 135
rect 227 133 229 135
rect 223 132 229 133
rect 236 132 240 134
rect 185 131 205 132
rect 173 128 174 130
rect 185 127 189 131
rect 236 130 237 132
rect 239 130 240 132
rect 280 134 300 135
rect 280 132 282 134
rect 284 132 300 134
rect 280 131 300 132
rect 177 123 189 127
rect 177 118 181 123
rect 177 116 178 118
rect 180 116 181 118
rect 177 104 181 116
rect 210 127 214 129
rect 210 125 211 127
rect 213 125 214 127
rect 210 119 214 125
rect 236 127 240 130
rect 236 123 260 127
rect 210 115 221 119
rect 177 101 194 104
rect 177 100 191 101
rect 190 99 191 100
rect 193 99 194 101
rect 179 96 185 97
rect 179 94 181 96
rect 183 94 185 96
rect 122 93 155 94
rect 122 91 151 93
rect 153 91 155 93
rect 122 90 155 91
rect 114 85 115 87
rect 117 85 118 87
rect 179 85 185 94
rect 190 94 194 99
rect 217 109 221 115
rect 256 119 260 123
rect 236 118 252 119
rect 236 116 248 118
rect 250 116 252 118
rect 236 115 252 116
rect 256 117 261 119
rect 256 115 258 117
rect 260 115 261 117
rect 236 109 240 115
rect 256 113 261 115
rect 256 111 260 113
rect 217 108 240 109
rect 217 106 219 108
rect 221 106 240 108
rect 217 105 240 106
rect 190 92 191 94
rect 193 92 194 94
rect 190 90 194 92
rect 199 94 205 95
rect 199 92 201 94
rect 203 92 205 94
rect 199 85 205 92
rect 228 94 232 96
rect 228 92 229 94
rect 231 92 232 94
rect 228 87 232 92
rect 236 94 240 105
rect 244 108 260 111
rect 244 106 245 108
rect 247 107 260 108
rect 296 127 300 131
rect 311 128 312 130
rect 296 123 308 127
rect 304 118 308 123
rect 304 116 305 118
rect 307 116 308 118
rect 247 106 248 107
rect 244 101 248 106
rect 244 99 245 101
rect 247 99 248 101
rect 244 97 248 99
rect 304 104 308 116
rect 291 101 308 104
rect 291 99 292 101
rect 294 100 308 101
rect 322 133 328 134
rect 322 131 324 133
rect 326 131 328 133
rect 322 130 328 131
rect 332 133 338 141
rect 332 131 334 133
rect 336 131 338 133
rect 349 135 364 136
rect 349 133 351 135
rect 353 133 364 135
rect 349 132 364 133
rect 332 130 338 131
rect 322 110 326 130
rect 360 127 364 132
rect 367 135 371 141
rect 367 133 368 135
rect 370 133 371 135
rect 367 131 371 133
rect 346 124 357 126
rect 346 122 354 124
rect 356 122 357 124
rect 360 125 374 127
rect 360 123 375 125
rect 346 120 357 122
rect 370 121 372 123
rect 374 121 375 123
rect 346 110 350 120
rect 370 119 375 121
rect 322 109 350 110
rect 322 107 324 109
rect 326 108 350 109
rect 326 107 347 108
rect 322 106 347 107
rect 349 106 350 108
rect 366 109 367 115
rect 346 104 350 106
rect 294 99 295 100
rect 280 94 286 95
rect 236 93 269 94
rect 236 91 265 93
rect 267 91 269 93
rect 236 90 269 91
rect 280 92 282 94
rect 284 92 286 94
rect 228 85 229 87
rect 231 85 232 87
rect 280 85 286 92
rect 291 94 295 99
rect 370 102 374 119
rect 358 98 374 102
rect 291 92 292 94
rect 294 92 295 94
rect 291 90 295 92
rect 300 96 306 97
rect 300 94 302 96
rect 304 94 306 96
rect 300 85 306 94
rect 349 97 362 98
rect 349 95 351 97
rect 353 95 362 97
rect 349 94 362 95
rect 400 135 404 141
rect 400 133 401 135
rect 403 133 404 135
rect 400 131 404 133
rect 407 135 422 136
rect 407 133 418 135
rect 420 133 422 135
rect 407 132 422 133
rect 433 133 439 141
rect 467 135 471 141
rect 407 127 411 132
rect 433 131 435 133
rect 437 131 439 133
rect 433 130 439 131
rect 443 133 449 134
rect 443 131 445 133
rect 447 131 449 133
rect 443 130 449 131
rect 397 125 411 127
rect 396 123 411 125
rect 414 124 425 126
rect 396 121 397 123
rect 399 121 401 123
rect 396 119 401 121
rect 414 122 415 124
rect 417 122 425 124
rect 414 120 425 122
rect 397 102 401 119
rect 404 109 405 115
rect 421 110 425 120
rect 445 110 449 130
rect 421 109 449 110
rect 421 108 445 109
rect 421 106 422 108
rect 424 107 445 108
rect 447 107 449 109
rect 424 106 449 107
rect 467 133 468 135
rect 470 133 471 135
rect 467 131 471 133
rect 474 135 489 136
rect 474 133 485 135
rect 487 133 489 135
rect 474 132 489 133
rect 500 133 506 141
rect 533 140 539 141
rect 533 138 535 140
rect 537 138 539 140
rect 533 137 539 138
rect 552 140 558 141
rect 552 138 554 140
rect 556 138 558 140
rect 552 137 558 138
rect 604 135 610 141
rect 474 127 478 132
rect 500 131 502 133
rect 504 131 506 133
rect 500 130 506 131
rect 510 133 516 134
rect 510 131 512 133
rect 514 131 516 133
rect 510 130 516 131
rect 464 125 478 127
rect 421 104 425 106
rect 397 98 413 102
rect 409 97 422 98
rect 409 95 418 97
rect 420 95 422 97
rect 409 94 422 95
rect 463 123 478 125
rect 481 124 492 126
rect 463 121 464 123
rect 466 121 468 123
rect 463 119 468 121
rect 481 122 482 124
rect 484 122 492 124
rect 481 120 492 122
rect 464 102 468 119
rect 471 109 472 115
rect 488 110 492 120
rect 512 110 516 130
rect 593 132 597 134
rect 604 133 606 135
rect 608 133 610 135
rect 604 132 610 133
rect 488 109 516 110
rect 488 108 512 109
rect 488 106 489 108
rect 491 107 512 108
rect 514 107 516 109
rect 491 106 516 107
rect 530 127 548 128
rect 530 125 544 127
rect 546 125 548 127
rect 530 124 548 125
rect 488 104 492 106
rect 530 118 534 124
rect 530 116 531 118
rect 533 116 534 118
rect 464 98 480 102
rect 476 97 489 98
rect 476 95 485 97
rect 487 95 489 97
rect 476 94 489 95
rect 526 95 527 106
rect 530 103 534 116
rect 593 130 594 132
rect 596 130 597 132
rect 593 127 597 130
rect 549 111 555 112
rect 530 99 545 103
rect 541 95 545 99
rect 573 123 597 127
rect 573 119 577 123
rect 619 127 623 129
rect 619 125 620 127
rect 622 125 623 127
rect 572 117 577 119
rect 572 115 573 117
rect 575 115 577 117
rect 581 118 597 119
rect 581 116 583 118
rect 585 116 597 118
rect 581 115 597 116
rect 572 113 577 115
rect 573 111 577 113
rect 573 108 589 111
rect 573 107 586 108
rect 585 106 586 107
rect 588 106 589 108
rect 585 101 589 106
rect 585 99 586 101
rect 588 99 589 101
rect 585 97 589 99
rect 593 109 597 115
rect 619 119 623 125
rect 612 115 623 119
rect 612 109 616 115
rect 593 108 616 109
rect 593 106 612 108
rect 614 106 616 108
rect 593 105 616 106
rect 541 94 558 95
rect 593 94 597 105
rect 541 92 554 94
rect 556 92 558 94
rect 541 91 558 92
rect 564 93 597 94
rect 564 91 566 93
rect 568 91 597 93
rect 564 90 597 91
rect 601 94 605 96
rect 601 92 602 94
rect 604 92 605 94
rect 333 87 337 89
rect 333 85 334 87
rect 336 85 337 87
rect 366 87 372 88
rect 366 85 368 87
rect 370 85 372 87
rect 399 87 405 88
rect 399 85 401 87
rect 403 85 405 87
rect 434 87 438 89
rect 434 85 435 87
rect 437 85 438 87
rect 466 87 472 88
rect 466 85 468 87
rect 470 85 472 87
rect 501 87 505 89
rect 501 85 502 87
rect 504 85 505 87
rect 533 87 539 88
rect 533 85 535 87
rect 537 85 539 87
rect 601 87 605 92
rect 601 85 602 87
rect 604 85 605 87
rect 17 67 19 69
rect 21 67 23 69
rect 17 66 23 67
rect 25 62 42 63
rect 25 60 38 62
rect 40 60 42 62
rect 25 59 42 60
rect 65 60 71 69
rect 10 48 11 59
rect 25 55 29 59
rect 65 58 67 60
rect 69 58 71 60
rect 65 57 71 58
rect 76 62 80 64
rect 76 60 77 62
rect 79 60 80 62
rect 14 51 29 55
rect 76 55 80 60
rect 85 62 91 69
rect 114 67 115 69
rect 117 67 118 69
rect 85 60 87 62
rect 89 60 91 62
rect 85 59 91 60
rect 114 62 118 67
rect 114 60 115 62
rect 117 60 118 62
rect 114 58 118 60
rect 122 63 155 64
rect 122 61 151 63
rect 153 61 155 63
rect 122 60 155 61
rect 179 60 185 69
rect 76 54 77 55
rect 14 38 18 51
rect 63 53 77 54
rect 79 53 80 55
rect 63 50 80 53
rect 33 42 39 43
rect 14 36 15 38
rect 17 36 18 38
rect 14 30 18 36
rect 14 29 32 30
rect 14 27 28 29
rect 30 27 32 29
rect 14 26 32 27
rect 63 38 67 50
rect 122 49 126 60
rect 179 58 181 60
rect 183 58 185 60
rect 179 57 185 58
rect 190 62 194 64
rect 190 60 191 62
rect 193 60 194 62
rect 103 48 126 49
rect 103 46 105 48
rect 107 46 126 48
rect 103 45 126 46
rect 103 39 107 45
rect 63 36 64 38
rect 66 36 67 38
rect 63 31 67 36
rect 63 27 75 31
rect 59 24 60 26
rect 71 23 75 27
rect 96 35 107 39
rect 96 29 100 35
rect 122 39 126 45
rect 130 55 134 57
rect 130 53 131 55
rect 133 53 134 55
rect 130 48 134 53
rect 130 46 131 48
rect 133 47 134 48
rect 133 46 146 47
rect 130 43 146 46
rect 142 41 146 43
rect 142 39 147 41
rect 122 38 138 39
rect 122 36 134 38
rect 136 36 138 38
rect 122 35 138 36
rect 142 37 144 39
rect 146 37 147 39
rect 142 35 147 37
rect 96 27 97 29
rect 99 27 100 29
rect 96 25 100 27
rect 142 31 146 35
rect 122 27 146 31
rect 122 24 126 27
rect 71 22 91 23
rect 122 22 123 24
rect 125 22 126 24
rect 71 20 87 22
rect 89 20 91 22
rect 71 19 91 20
rect 109 21 115 22
rect 109 19 111 21
rect 113 19 115 21
rect 122 20 126 22
rect 190 55 194 60
rect 199 62 205 69
rect 228 67 229 69
rect 231 67 232 69
rect 199 60 201 62
rect 203 60 205 62
rect 199 59 205 60
rect 228 62 232 67
rect 228 60 229 62
rect 231 60 232 62
rect 228 58 232 60
rect 236 63 269 64
rect 236 61 265 63
rect 267 61 269 63
rect 236 60 269 61
rect 280 62 286 69
rect 280 60 282 62
rect 284 60 286 62
rect 190 54 191 55
rect 177 53 191 54
rect 193 53 194 55
rect 177 50 194 53
rect 177 38 181 50
rect 236 49 240 60
rect 280 59 286 60
rect 291 62 295 64
rect 291 60 292 62
rect 294 60 295 62
rect 217 48 240 49
rect 217 46 219 48
rect 221 46 240 48
rect 217 45 240 46
rect 217 39 221 45
rect 177 36 178 38
rect 180 36 181 38
rect 177 31 181 36
rect 177 27 189 31
rect 173 24 174 26
rect 17 16 23 17
rect 17 14 19 16
rect 21 14 23 16
rect 17 13 23 14
rect 36 16 42 17
rect 36 14 38 16
rect 40 14 42 16
rect 36 13 42 14
rect 109 13 115 19
rect 185 23 189 27
rect 210 35 221 39
rect 210 29 214 35
rect 236 39 240 45
rect 244 55 248 57
rect 244 53 245 55
rect 247 53 248 55
rect 244 48 248 53
rect 244 46 245 48
rect 247 47 248 48
rect 247 46 260 47
rect 244 43 260 46
rect 256 41 260 43
rect 291 55 295 60
rect 300 60 306 69
rect 333 67 334 69
rect 336 67 337 69
rect 333 65 337 67
rect 366 67 368 69
rect 370 67 372 69
rect 366 66 372 67
rect 399 67 401 69
rect 403 67 405 69
rect 399 66 405 67
rect 434 67 435 69
rect 437 67 438 69
rect 434 65 438 67
rect 466 67 468 69
rect 470 67 472 69
rect 466 66 472 67
rect 501 67 502 69
rect 504 67 505 69
rect 501 65 505 67
rect 533 67 535 69
rect 537 67 539 69
rect 533 66 539 67
rect 601 67 602 69
rect 604 67 605 69
rect 300 58 302 60
rect 304 58 306 60
rect 300 57 306 58
rect 291 53 292 55
rect 294 54 295 55
rect 294 53 308 54
rect 291 50 308 53
rect 256 39 261 41
rect 236 38 252 39
rect 236 36 248 38
rect 250 36 252 38
rect 236 35 252 36
rect 256 37 258 39
rect 260 37 261 39
rect 256 35 261 37
rect 210 27 211 29
rect 213 27 214 29
rect 210 25 214 27
rect 256 31 260 35
rect 236 27 260 31
rect 236 24 240 27
rect 185 22 205 23
rect 236 22 237 24
rect 239 22 240 24
rect 304 38 308 50
rect 349 59 362 60
rect 349 57 351 59
rect 353 57 362 59
rect 349 56 362 57
rect 358 52 374 56
rect 346 48 350 50
rect 304 36 305 38
rect 307 36 308 38
rect 304 31 308 36
rect 296 27 308 31
rect 296 23 300 27
rect 311 24 312 26
rect 185 20 201 22
rect 203 20 205 22
rect 185 19 205 20
rect 223 21 229 22
rect 223 19 225 21
rect 227 19 229 21
rect 236 20 240 22
rect 280 22 300 23
rect 280 20 282 22
rect 284 20 300 22
rect 280 19 300 20
rect 223 13 229 19
rect 322 47 347 48
rect 322 45 324 47
rect 326 46 347 47
rect 349 46 350 48
rect 326 45 350 46
rect 322 44 350 45
rect 322 24 326 44
rect 346 34 350 44
rect 366 39 367 45
rect 370 35 374 52
rect 346 32 357 34
rect 346 30 354 32
rect 356 30 357 32
rect 370 33 375 35
rect 370 31 372 33
rect 374 31 375 33
rect 346 28 357 30
rect 360 29 375 31
rect 360 27 374 29
rect 322 23 328 24
rect 322 21 324 23
rect 326 21 328 23
rect 322 20 328 21
rect 332 23 338 24
rect 332 21 334 23
rect 336 21 338 23
rect 360 22 364 27
rect 332 13 338 21
rect 349 21 364 22
rect 349 19 351 21
rect 353 19 364 21
rect 349 18 364 19
rect 367 21 371 23
rect 367 19 368 21
rect 370 19 371 21
rect 367 13 371 19
rect 409 59 422 60
rect 409 57 418 59
rect 420 57 422 59
rect 409 56 422 57
rect 397 52 413 56
rect 397 35 401 52
rect 476 59 489 60
rect 421 48 425 50
rect 404 39 405 45
rect 421 46 422 48
rect 424 47 449 48
rect 424 46 445 47
rect 421 45 445 46
rect 447 45 449 47
rect 421 44 449 45
rect 396 33 401 35
rect 421 34 425 44
rect 396 31 397 33
rect 399 31 401 33
rect 414 32 425 34
rect 396 29 411 31
rect 397 27 411 29
rect 414 30 415 32
rect 417 30 425 32
rect 414 28 425 30
rect 400 21 404 23
rect 400 19 401 21
rect 403 19 404 21
rect 400 13 404 19
rect 407 22 411 27
rect 445 24 449 44
rect 433 23 439 24
rect 407 21 422 22
rect 407 19 418 21
rect 420 19 422 21
rect 407 18 422 19
rect 433 21 435 23
rect 437 21 439 23
rect 433 13 439 21
rect 443 23 449 24
rect 443 21 445 23
rect 447 21 449 23
rect 443 20 449 21
rect 476 57 485 59
rect 487 57 489 59
rect 476 56 489 57
rect 464 52 480 56
rect 464 35 468 52
rect 564 63 597 64
rect 541 62 558 63
rect 541 60 554 62
rect 556 60 558 62
rect 564 61 566 63
rect 568 61 597 63
rect 564 60 597 61
rect 541 59 558 60
rect 488 48 492 50
rect 471 39 472 45
rect 488 46 489 48
rect 491 47 516 48
rect 491 46 512 47
rect 488 45 512 46
rect 514 45 516 47
rect 488 44 516 45
rect 463 33 468 35
rect 488 34 492 44
rect 463 31 464 33
rect 466 31 468 33
rect 481 32 492 34
rect 463 29 478 31
rect 464 27 478 29
rect 481 30 482 32
rect 484 30 492 32
rect 481 28 492 30
rect 467 21 471 23
rect 467 19 468 21
rect 470 19 471 21
rect 467 13 471 19
rect 474 22 478 27
rect 512 24 516 44
rect 526 48 527 59
rect 541 55 545 59
rect 530 51 545 55
rect 530 38 534 51
rect 585 55 589 57
rect 585 53 586 55
rect 588 53 589 55
rect 549 42 555 43
rect 530 36 531 38
rect 533 36 534 38
rect 530 30 534 36
rect 530 29 548 30
rect 530 27 544 29
rect 546 27 548 29
rect 530 26 548 27
rect 585 48 589 53
rect 585 47 586 48
rect 573 46 586 47
rect 588 46 589 48
rect 573 43 589 46
rect 593 49 597 60
rect 601 62 605 67
rect 601 60 602 62
rect 604 60 605 62
rect 601 58 605 60
rect 593 48 616 49
rect 593 46 612 48
rect 614 46 616 48
rect 593 45 616 46
rect 573 41 577 43
rect 572 39 577 41
rect 593 39 597 45
rect 572 37 573 39
rect 575 37 577 39
rect 572 35 577 37
rect 581 38 597 39
rect 581 36 583 38
rect 585 36 597 38
rect 581 35 597 36
rect 500 23 506 24
rect 474 21 489 22
rect 474 19 485 21
rect 487 19 489 21
rect 474 18 489 19
rect 500 21 502 23
rect 504 21 506 23
rect 500 13 506 21
rect 510 23 516 24
rect 510 21 512 23
rect 514 21 516 23
rect 510 20 516 21
rect 573 31 577 35
rect 612 39 616 45
rect 612 35 623 39
rect 573 27 597 31
rect 593 24 597 27
rect 619 29 623 35
rect 619 27 620 29
rect 622 27 623 29
rect 619 25 623 27
rect 593 22 594 24
rect 596 22 597 24
rect 593 20 597 22
rect 604 21 610 22
rect 604 19 606 21
rect 608 19 610 21
rect 533 16 539 17
rect 533 14 535 16
rect 537 14 539 16
rect 533 13 539 14
rect 552 16 558 17
rect 552 14 554 16
rect 556 14 558 16
rect 552 13 558 14
rect 604 13 610 19
<< via1 >>
rect 39 548 41 550
rect 80 557 82 559
rect 105 557 107 559
rect 88 533 90 535
rect 152 556 154 558
rect 97 533 99 535
rect 170 548 172 550
rect 194 557 196 559
rect 219 557 221 559
rect 202 533 204 535
rect 211 533 213 535
rect 266 541 268 543
rect 313 556 315 558
rect 330 556 332 558
rect 355 540 357 542
rect 332 532 334 534
rect 379 548 381 550
rect 406 548 408 550
rect 437 556 439 558
rect 457 556 459 558
rect 480 541 482 543
rect 505 556 507 558
rect 523 540 525 542
rect 504 532 506 534
rect 565 556 567 558
rect 88 483 90 485
rect 39 468 41 470
rect 97 483 99 485
rect 80 459 82 461
rect 105 459 107 461
rect 152 460 154 462
rect 202 483 204 485
rect 170 468 172 470
rect 211 483 213 485
rect 194 459 196 461
rect 266 475 268 477
rect 219 459 221 461
rect 332 484 334 486
rect 313 460 315 462
rect 330 460 332 462
rect 355 476 357 478
rect 379 468 381 470
rect 406 468 408 470
rect 437 460 439 462
rect 504 484 506 486
rect 480 475 482 477
rect 457 460 459 462
rect 505 460 507 462
rect 523 476 525 478
rect 565 460 567 462
rect 39 404 41 406
rect 80 413 82 415
rect 105 413 107 415
rect 88 389 90 391
rect 152 412 154 414
rect 97 389 99 391
rect 170 404 172 406
rect 194 413 196 415
rect 219 413 221 415
rect 202 389 204 391
rect 211 389 213 391
rect 266 397 268 399
rect 313 412 315 414
rect 330 412 332 414
rect 355 396 357 398
rect 332 388 334 390
rect 379 404 381 406
rect 406 404 408 406
rect 437 412 439 414
rect 457 412 459 414
rect 480 397 482 399
rect 505 412 507 414
rect 523 396 525 398
rect 504 388 506 390
rect 565 412 567 414
rect 88 339 90 341
rect 39 324 41 326
rect 97 339 99 341
rect 80 315 82 317
rect 105 315 107 317
rect 152 316 154 318
rect 202 339 204 341
rect 170 324 172 326
rect 211 339 213 341
rect 194 315 196 317
rect 266 331 268 333
rect 219 315 221 317
rect 332 340 334 342
rect 313 316 315 318
rect 330 316 332 318
rect 355 332 357 334
rect 379 324 381 326
rect 406 324 408 326
rect 437 316 439 318
rect 504 340 506 342
rect 480 331 482 333
rect 457 316 459 318
rect 505 316 507 318
rect 523 332 525 334
rect 565 316 567 318
rect 39 260 41 262
rect 80 269 82 271
rect 105 269 107 271
rect 88 245 90 247
rect 152 268 154 270
rect 97 245 99 247
rect 170 260 172 262
rect 194 269 196 271
rect 219 269 221 271
rect 202 245 204 247
rect 211 245 213 247
rect 266 253 268 255
rect 313 268 315 270
rect 330 268 332 270
rect 355 252 357 254
rect 332 244 334 246
rect 379 260 381 262
rect 406 260 408 262
rect 437 268 439 270
rect 457 268 459 270
rect 480 253 482 255
rect 505 268 507 270
rect 523 252 525 254
rect 504 244 506 246
rect 565 268 567 270
rect 88 195 90 197
rect 39 180 41 182
rect 97 195 99 197
rect 80 171 82 173
rect 105 171 107 173
rect 152 172 154 174
rect 202 195 204 197
rect 170 180 172 182
rect 211 195 213 197
rect 194 171 196 173
rect 266 187 268 189
rect 219 171 221 173
rect 332 196 334 198
rect 313 172 315 174
rect 330 172 332 174
rect 355 188 357 190
rect 379 180 381 182
rect 406 180 408 182
rect 437 172 439 174
rect 504 196 506 198
rect 480 187 482 189
rect 457 172 459 174
rect 505 172 507 174
rect 523 188 525 190
rect 565 172 567 174
rect 39 116 41 118
rect 80 125 82 127
rect 105 125 107 127
rect 88 101 90 103
rect 152 124 154 126
rect 97 101 99 103
rect 170 116 172 118
rect 194 125 196 127
rect 219 125 221 127
rect 202 101 204 103
rect 211 101 213 103
rect 266 109 268 111
rect 313 124 315 126
rect 330 124 332 126
rect 355 108 357 110
rect 332 100 334 102
rect 379 116 381 118
rect 406 116 408 118
rect 437 124 439 126
rect 457 124 459 126
rect 480 109 482 111
rect 505 124 507 126
rect 523 108 525 110
rect 504 100 506 102
rect 565 124 567 126
rect 88 51 90 53
rect 39 36 41 38
rect 97 51 99 53
rect 80 27 82 29
rect 105 27 107 29
rect 152 28 154 30
rect 202 51 204 53
rect 170 36 172 38
rect 211 51 213 53
rect 194 27 196 29
rect 266 43 268 45
rect 219 27 221 29
rect 332 52 334 54
rect 313 28 315 30
rect 330 28 332 30
rect 355 44 357 46
rect 379 36 381 38
rect 406 36 408 38
rect 437 28 439 30
rect 504 52 506 54
rect 480 43 482 45
rect 457 28 459 30
rect 505 28 507 30
rect 523 44 525 46
rect 565 28 567 30
<< labels >>
rlabel alu1 125 9 125 9 6 vss
rlabel alu1 125 73 125 73 6 vdd
rlabel alu1 73 73 73 73 6 vdd
rlabel alu1 73 9 73 9 6 vss
rlabel alu1 239 9 239 9 6 vss
rlabel alu1 239 73 239 73 6 vdd
rlabel alu1 187 73 187 73 6 vdd
rlabel alu1 187 9 187 9 6 vss
rlabel alu1 24 9 24 9 6 vss
rlabel alu1 24 73 24 73 6 vdd
rlabel via1 204 52 204 52 1 cin
rlabel alu1 298 9 298 9 4 vss
rlabel alu1 298 73 298 73 4 vdd
rlabel alu1 419 9 419 9 6 vss
rlabel alu1 419 73 419 73 6 vdd
rlabel alu1 352 9 352 9 4 vss
rlabel alu1 352 73 352 73 4 vdd
rlabel alu1 486 9 486 9 6 vss
rlabel alu1 486 73 486 73 6 vdd
rlabel via1 506 53 506 53 1 s1
rlabel alu1 514 61 514 61 1 s1
rlabel via1 332 53 332 53 1 s1
rlabel alu1 324 61 324 61 1 s1
rlabel alu1 447 61 447 61 1 s0
rlabel alu1 540 9 540 9 6 vss
rlabel alu1 540 73 540 73 6 vdd
rlabel alu1 594 9 594 9 4 vss
rlabel alu1 594 73 594 73 4 vdd
rlabel alu1 80 33 80 33 1 a0
rlabel via1 88 51 88 51 1 b0
rlabel alu1 282 53 282 53 1 b0
rlabel alu1 298 37 298 37 1 a0
rlabel alu1 540 37 540 37 1 a0
rlabel alu1 548 37 548 37 1 a0
rlabel alu1 540 45 540 45 1 b0
rlabel alu1 548 45 548 45 1 b0
rlabel alu1 556 53 556 53 1 b0
rlabel alu1 614 61 614 61 1 b0
rlabel alu1 622 53 622 53 1 b0
rlabel polyct1 606 33 606 33 1 a0
rlabel alu1 614 29 614 29 1 a0
rlabel alu1 290 33 290 33 1 a0
rlabel alu1 391 47 391 47 1 z0
rlabel alu1 399 61 399 61 1 z0
rlabel alu1 125 145 125 145 8 vss
rlabel alu1 125 81 125 81 8 vdd
rlabel alu1 73 81 73 81 8 vdd
rlabel alu1 73 145 73 145 8 vss
rlabel alu1 239 145 239 145 8 vss
rlabel alu1 239 81 239 81 8 vdd
rlabel alu1 187 81 187 81 8 vdd
rlabel alu1 187 145 187 145 8 vss
rlabel alu1 24 145 24 145 8 vss
rlabel alu1 24 81 24 81 8 vdd
rlabel alu1 298 145 298 145 2 vss
rlabel alu1 298 81 298 81 2 vdd
rlabel alu1 419 145 419 145 8 vss
rlabel alu1 419 81 419 81 8 vdd
rlabel alu1 352 145 352 145 2 vss
rlabel alu1 352 81 352 81 2 vdd
rlabel alu1 486 145 486 145 8 vss
rlabel alu1 486 81 486 81 8 vdd
rlabel via1 506 101 506 101 5 s1
rlabel alu1 514 93 514 93 5 s1
rlabel via1 332 101 332 101 5 s1
rlabel alu1 324 93 324 93 5 s1
rlabel alu1 447 93 447 93 5 s0
rlabel alu1 540 145 540 145 8 vss
rlabel alu1 540 81 540 81 8 vdd
rlabel alu1 594 145 594 145 2 vss
rlabel alu1 594 81 594 81 2 vdd
rlabel via1 204 102 204 102 1 cin1
rlabel alu1 8 39 8 39 1 cin1
rlabel alu1 80 121 80 121 1 a1
rlabel via1 88 103 88 103 1 b1
rlabel alu1 282 101 282 101 1 b1
rlabel alu1 290 121 290 121 1 a1
rlabel alu1 298 117 298 117 1 a1
rlabel alu1 391 107 391 107 1 z1
rlabel alu1 399 93 399 93 1 z1
rlabel alu1 540 117 540 117 1 a1
rlabel alu1 548 117 548 117 1 a1
rlabel alu1 540 109 540 109 1 b1
rlabel alu1 548 109 548 109 1 b1
rlabel alu1 556 101 556 101 1 b1
rlabel polyct1 606 121 606 121 1 a1
rlabel alu1 614 125 614 125 1 a1
rlabel alu1 622 101 622 101 1 b1
rlabel alu1 614 93 614 93 1 b1
rlabel alu1 8 115 8 115 1 cin2
rlabel alu1 125 153 125 153 6 vss
rlabel alu1 125 217 125 217 6 vdd
rlabel alu1 73 217 73 217 6 vdd
rlabel alu1 73 153 73 153 6 vss
rlabel alu1 239 153 239 153 6 vss
rlabel alu1 239 217 239 217 6 vdd
rlabel alu1 187 217 187 217 6 vdd
rlabel alu1 187 153 187 153 6 vss
rlabel alu1 24 153 24 153 6 vss
rlabel alu1 24 217 24 217 6 vdd
rlabel alu1 298 153 298 153 4 vss
rlabel alu1 298 217 298 217 4 vdd
rlabel alu1 419 153 419 153 6 vss
rlabel alu1 419 217 419 217 6 vdd
rlabel alu1 352 153 352 153 4 vss
rlabel alu1 352 217 352 217 4 vdd
rlabel alu1 486 153 486 153 6 vss
rlabel alu1 486 217 486 217 6 vdd
rlabel via1 506 197 506 197 1 s1
rlabel alu1 514 205 514 205 1 s1
rlabel via1 332 197 332 197 1 s1
rlabel alu1 324 205 324 205 1 s1
rlabel alu1 447 205 447 205 1 s0
rlabel alu1 540 153 540 153 6 vss
rlabel alu1 540 217 540 217 6 vdd
rlabel alu1 594 153 594 153 4 vss
rlabel alu1 594 217 594 217 4 vdd
rlabel alu1 125 225 125 225 8 vdd
rlabel alu1 73 225 73 225 8 vdd
rlabel alu1 239 225 239 225 8 vdd
rlabel alu1 187 225 187 225 8 vdd
rlabel alu1 24 225 24 225 8 vdd
rlabel alu1 298 225 298 225 2 vdd
rlabel alu1 419 225 419 225 8 vdd
rlabel alu1 352 225 352 225 2 vdd
rlabel alu1 486 225 486 225 8 vdd
rlabel via1 506 245 506 245 5 s1
rlabel alu1 514 237 514 237 5 s1
rlabel via1 332 245 332 245 5 s1
rlabel alu1 324 237 324 237 5 s1
rlabel alu1 447 237 447 237 5 s0
rlabel alu1 540 225 540 225 8 vdd
rlabel alu1 594 225 594 225 2 vdd
rlabel alu1 8 183 8 183 1 cin3
rlabel alu1 80 177 80 177 1 a2
rlabel via1 88 195 88 195 1 b2
rlabel alu1 282 197 282 197 1 b2
rlabel alu1 290 177 290 177 1 a2
rlabel alu1 298 181 298 181 1 a2
rlabel alu1 391 191 391 191 1 z2
rlabel alu1 399 205 399 205 1 z2
rlabel alu1 540 181 540 181 1 a2
rlabel alu1 548 181 548 181 1 a2
rlabel alu1 540 189 540 189 1 b2
rlabel alu1 548 189 548 189 1 b2
rlabel alu1 556 197 556 197 1 b2
rlabel alu1 614 205 614 205 1 b2
rlabel alu1 622 197 622 197 1 b2
rlabel polyct1 606 177 606 177 1 a2
rlabel alu1 614 173 614 173 1 a2
rlabel via1 204 196 204 196 1 cin2
rlabel via1 88 247 88 247 1 b3
rlabel alu1 80 265 80 265 1 a3
rlabel via1 204 246 204 246 1 cin3
rlabel alu1 282 245 282 245 1 b3
rlabel alu1 290 265 290 265 1 a3
rlabel alu1 298 261 298 261 1 a3
rlabel alu1 391 251 391 251 1 z3
rlabel alu1 399 237 399 237 1 z3
rlabel alu1 540 261 540 261 1 a3
rlabel alu1 548 261 548 261 1 a3
rlabel alu1 540 253 540 253 1 b3
rlabel alu1 548 253 548 253 1 b3
rlabel alu1 556 245 556 245 1 b3
rlabel polyct1 606 265 606 265 1 a3
rlabel alu1 614 237 614 237 1 b3
rlabel alu1 622 245 622 245 1 b3
rlabel alu1 8 259 8 259 1 cin4
rlabel alu1 614 269 614 269 1 a3
rlabel alu1 594 289 594 289 2 vss
rlabel alu1 540 289 540 289 8 vss
rlabel alu1 486 289 486 289 8 vss
rlabel alu1 352 289 352 289 2 vss
rlabel alu1 419 289 419 289 8 vss
rlabel alu1 298 289 298 289 2 vss
rlabel alu1 24 289 24 289 8 vss
rlabel alu1 187 289 187 289 8 vss
rlabel alu1 239 289 239 289 8 vss
rlabel alu1 73 289 73 289 8 vss
rlabel alu1 125 289 125 289 8 vss
rlabel alu1 125 297 125 297 6 vss
rlabel alu1 125 361 125 361 6 vdd
rlabel alu1 73 361 73 361 6 vdd
rlabel alu1 73 297 73 297 6 vss
rlabel alu1 239 297 239 297 6 vss
rlabel alu1 239 361 239 361 6 vdd
rlabel alu1 187 361 187 361 6 vdd
rlabel alu1 187 297 187 297 6 vss
rlabel alu1 24 297 24 297 6 vss
rlabel alu1 24 361 24 361 6 vdd
rlabel alu1 298 297 298 297 4 vss
rlabel alu1 298 361 298 361 4 vdd
rlabel alu1 419 297 419 297 6 vss
rlabel alu1 419 361 419 361 6 vdd
rlabel alu1 352 297 352 297 4 vss
rlabel alu1 352 361 352 361 4 vdd
rlabel alu1 486 297 486 297 6 vss
rlabel alu1 486 361 486 361 6 vdd
rlabel via1 506 341 506 341 1 s1
rlabel alu1 514 349 514 349 1 s1
rlabel via1 332 341 332 341 1 s1
rlabel alu1 324 349 324 349 1 s1
rlabel alu1 447 349 447 349 1 s0
rlabel alu1 540 297 540 297 6 vss
rlabel alu1 540 361 540 361 6 vdd
rlabel alu1 594 297 594 297 4 vss
rlabel alu1 594 361 594 361 4 vdd
rlabel alu1 125 433 125 433 8 vss
rlabel alu1 125 369 125 369 8 vdd
rlabel alu1 73 369 73 369 8 vdd
rlabel alu1 73 433 73 433 8 vss
rlabel alu1 239 433 239 433 8 vss
rlabel alu1 239 369 239 369 8 vdd
rlabel alu1 187 369 187 369 8 vdd
rlabel alu1 187 433 187 433 8 vss
rlabel alu1 24 433 24 433 8 vss
rlabel alu1 24 369 24 369 8 vdd
rlabel alu1 298 433 298 433 2 vss
rlabel alu1 298 369 298 369 2 vdd
rlabel alu1 419 433 419 433 8 vss
rlabel alu1 419 369 419 369 8 vdd
rlabel alu1 352 433 352 433 2 vss
rlabel alu1 352 369 352 369 2 vdd
rlabel alu1 486 433 486 433 8 vss
rlabel alu1 486 369 486 369 8 vdd
rlabel via1 506 389 506 389 5 s1
rlabel alu1 514 381 514 381 5 s1
rlabel via1 332 389 332 389 5 s1
rlabel alu1 324 381 324 381 5 s1
rlabel alu1 447 381 447 381 5 s0
rlabel alu1 540 433 540 433 8 vss
rlabel alu1 540 369 540 369 8 vdd
rlabel alu1 594 433 594 433 2 vss
rlabel alu1 594 369 594 369 2 vdd
rlabel alu1 125 441 125 441 6 vss
rlabel alu1 125 505 125 505 6 vdd
rlabel alu1 73 505 73 505 6 vdd
rlabel alu1 73 441 73 441 6 vss
rlabel alu1 239 441 239 441 6 vss
rlabel alu1 239 505 239 505 6 vdd
rlabel alu1 187 505 187 505 6 vdd
rlabel alu1 187 441 187 441 6 vss
rlabel alu1 24 441 24 441 6 vss
rlabel alu1 24 505 24 505 6 vdd
rlabel alu1 298 441 298 441 4 vss
rlabel alu1 298 505 298 505 4 vdd
rlabel alu1 419 441 419 441 6 vss
rlabel alu1 419 505 419 505 6 vdd
rlabel alu1 352 441 352 441 4 vss
rlabel alu1 352 505 352 505 4 vdd
rlabel alu1 486 441 486 441 6 vss
rlabel alu1 486 505 486 505 6 vdd
rlabel via1 506 485 506 485 1 s1
rlabel alu1 514 493 514 493 1 s1
rlabel via1 332 485 332 485 1 s1
rlabel alu1 324 493 324 493 1 s1
rlabel alu1 447 493 447 493 1 s0
rlabel alu1 540 441 540 441 6 vss
rlabel alu1 540 505 540 505 6 vdd
rlabel alu1 594 441 594 441 4 vss
rlabel alu1 594 505 594 505 4 vdd
rlabel alu1 125 577 125 577 8 vss
rlabel alu1 125 513 125 513 8 vdd
rlabel alu1 73 513 73 513 8 vdd
rlabel alu1 73 577 73 577 8 vss
rlabel alu1 239 577 239 577 8 vss
rlabel alu1 239 513 239 513 8 vdd
rlabel alu1 187 513 187 513 8 vdd
rlabel alu1 187 577 187 577 8 vss
rlabel alu1 24 577 24 577 8 vss
rlabel alu1 24 513 24 513 8 vdd
rlabel alu1 8 547 8 547 5 cout
rlabel alu1 298 577 298 577 2 vss
rlabel alu1 298 513 298 513 2 vdd
rlabel alu1 419 577 419 577 8 vss
rlabel alu1 419 513 419 513 8 vdd
rlabel alu1 352 577 352 577 2 vss
rlabel alu1 352 513 352 513 2 vdd
rlabel alu1 486 577 486 577 8 vss
rlabel alu1 486 513 486 513 8 vdd
rlabel via1 506 533 506 533 5 s1
rlabel alu1 514 525 514 525 5 s1
rlabel via1 332 533 332 533 5 s1
rlabel alu1 324 525 324 525 5 s1
rlabel alu1 447 525 447 525 5 s0
rlabel alu1 540 577 540 577 8 vss
rlabel alu1 540 513 540 513 8 vdd
rlabel alu1 594 577 594 577 2 vss
rlabel alu1 594 513 594 513 2 vdd
rlabel alu1 80 321 80 321 1 a4
rlabel via1 88 339 88 339 1 b4
rlabel alu1 8 327 8 327 1 cin5
rlabel via1 204 340 204 340 1 cin4
rlabel alu1 282 341 282 341 1 b4
rlabel alu1 290 321 290 321 1 a4
rlabel alu1 298 325 298 325 1 a4
rlabel alu1 391 335 391 335 1 z4
rlabel alu1 399 349 399 349 1 z4
rlabel alu1 540 333 540 333 1 b4
rlabel alu1 548 333 548 333 1 b4
rlabel alu1 556 341 556 341 1 b4
rlabel alu1 540 325 540 325 1 a4
rlabel alu1 548 325 548 325 1 a4
rlabel polyct1 606 321 606 321 1 a4
rlabel alu1 614 317 614 317 1 a4
rlabel alu1 614 349 614 349 1 b4
rlabel alu1 622 341 622 341 1 b4
rlabel alu1 614 381 614 381 1 b5
rlabel alu1 622 389 622 389 1 b5
rlabel polyct1 606 409 606 409 1 a5
rlabel alu1 614 413 614 413 1 a5
rlabel alu1 540 405 540 405 1 a5
rlabel alu1 548 405 548 405 1 a5
rlabel alu1 540 397 540 397 1 b5
rlabel alu1 548 397 548 397 1 b5
rlabel alu1 556 389 556 389 1 b5
rlabel alu1 391 395 391 395 1 z5
rlabel alu1 399 381 399 381 1 z5
rlabel alu1 290 409 290 409 1 a5
rlabel alu1 298 405 298 405 1 a5
rlabel alu1 282 389 282 389 1 b5
rlabel via1 204 390 204 390 1 cin5
rlabel alu1 80 409 80 409 1 a5
rlabel via1 88 391 88 391 1 b5
rlabel alu1 8 403 8 403 1 cin6
rlabel alu1 80 465 80 465 1 a6
rlabel via1 88 483 88 483 1 b6
rlabel via1 204 484 204 484 1 cin6
rlabel alu1 282 485 282 485 1 b6
rlabel alu1 290 465 290 465 1 a6
rlabel alu1 298 469 298 469 1 a6
rlabel alu1 391 479 391 479 1 z6
rlabel alu1 399 493 399 493 1 z6
rlabel alu1 540 469 540 469 1 a6
rlabel alu1 548 469 548 469 1 a6
rlabel alu1 540 477 540 477 1 b6
rlabel alu1 548 477 548 477 1 b6
rlabel alu1 556 485 556 485 1 b6
rlabel polyct1 606 465 606 465 1 a6
rlabel alu1 614 461 614 461 1 a6
rlabel alu1 614 493 614 493 1 b6
rlabel alu1 622 485 622 485 1 b6
rlabel alu1 80 553 80 553 1 a7
rlabel via1 88 535 88 535 1 b7
rlabel alu1 8 471 8 471 1 cin7
rlabel via1 204 534 204 534 1 cin7
rlabel alu1 282 533 282 533 1 b7
rlabel alu1 290 553 290 553 1 a7
rlabel alu1 298 549 298 549 1 a7
rlabel alu1 540 549 540 549 1 a7
rlabel alu1 548 549 548 549 1 a7
rlabel polyct1 606 553 606 553 1 a7
rlabel alu1 614 557 614 557 1 a7
rlabel alu1 540 541 540 541 1 b7
rlabel alu1 548 541 548 541 1 b7
rlabel alu1 556 533 556 533 1 b7
rlabel alu1 614 525 614 525 1 b7
rlabel alu1 622 533 622 533 1 b7
rlabel alu1 391 539 391 539 1 z7
rlabel alu1 399 525 399 525 1 z7
<< end >>
