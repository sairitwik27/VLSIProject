magic
tech scmos
timestamp 1608918681
<< ab >>
rect 9 141 57 149
rect 18 76 57 141
rect 59 76 95 149
rect 18 13 55 76
rect 9 5 55 13
rect 57 5 95 76
rect 97 141 102 149
rect 97 85 99 141
rect 97 76 102 85
rect 104 76 167 149
rect 169 141 262 149
rect 169 117 207 141
rect 169 85 216 117
rect 223 85 262 141
rect 169 76 262 85
rect 264 76 300 149
rect 97 5 137 76
rect 139 5 202 76
rect 207 69 260 76
rect 207 37 216 69
rect 223 13 260 69
rect 204 5 260 13
rect 262 5 300 76
rect 302 141 307 149
rect 302 85 304 141
rect 302 76 307 85
rect 309 76 372 149
rect 374 117 412 149
rect 374 76 421 117
rect 302 5 342 76
rect 344 5 407 76
rect 412 37 421 76
rect -249 -67 -169 5
rect -167 -67 -64 5
rect -62 -67 81 5
rect 83 -67 186 5
rect 188 -67 331 5
rect 333 -67 436 5
rect 438 -67 581 5
rect 583 -67 686 5
rect 688 -67 751 5
<< nwell >>
rect 0 37 421 117
rect -254 -72 756 -27
<< pwell >>
rect 0 117 421 154
rect 0 10 421 37
rect -254 -27 756 10
<< poly >>
rect 26 136 28 141
rect 33 136 35 141
rect 46 134 48 138
rect 66 136 68 141
rect 73 136 75 141
rect 131 145 156 147
rect 114 140 116 145
rect 121 140 123 145
rect 86 134 88 138
rect 131 137 133 145
rect 141 137 143 141
rect 154 137 156 145
rect 154 135 159 137
rect 178 136 180 141
rect 185 136 187 141
rect 157 132 159 135
rect 26 112 28 125
rect 33 120 35 125
rect 46 120 48 125
rect 32 118 38 120
rect 32 116 34 118
rect 36 116 38 118
rect 32 114 38 116
rect 42 118 48 120
rect 42 116 44 118
rect 46 116 48 118
rect 42 114 48 116
rect 22 110 28 112
rect 22 108 24 110
rect 26 108 28 110
rect 22 106 28 108
rect 26 103 28 106
rect 36 103 38 114
rect 46 110 48 114
rect 66 112 68 125
rect 73 120 75 125
rect 86 120 88 125
rect 72 118 78 120
rect 72 116 74 118
rect 76 116 78 118
rect 72 114 78 116
rect 82 118 88 120
rect 114 119 116 128
rect 121 125 123 128
rect 121 123 125 125
rect 131 124 133 128
rect 141 125 143 128
rect 123 120 125 123
rect 141 123 150 125
rect 198 134 200 138
rect 231 136 233 141
rect 238 136 240 141
rect 251 134 253 138
rect 271 136 273 141
rect 278 136 280 141
rect 336 145 361 147
rect 319 140 321 145
rect 326 140 328 145
rect 291 134 293 138
rect 336 137 338 145
rect 346 137 348 141
rect 359 137 361 145
rect 359 135 364 137
rect 383 136 385 141
rect 390 136 392 141
rect 362 132 364 135
rect 141 121 146 123
rect 148 121 150 123
rect 82 116 84 118
rect 86 116 88 118
rect 82 114 88 116
rect 62 110 68 112
rect 62 108 64 110
rect 66 108 68 110
rect 62 106 68 108
rect 66 103 68 106
rect 76 103 78 114
rect 86 110 88 114
rect 113 117 119 119
rect 113 115 115 117
rect 117 115 119 117
rect 113 113 119 115
rect 123 118 129 120
rect 123 116 125 118
rect 127 116 129 118
rect 123 114 129 116
rect 141 119 150 121
rect 141 115 143 119
rect 157 115 159 123
rect 113 110 115 113
rect 123 110 125 114
rect 133 113 143 115
rect 149 113 162 115
rect 133 110 135 113
rect 149 110 151 113
rect 160 112 162 113
rect 178 112 180 125
rect 185 120 187 125
rect 198 120 200 125
rect 184 118 190 120
rect 184 116 186 118
rect 188 116 190 118
rect 184 114 190 116
rect 194 118 200 120
rect 194 116 196 118
rect 198 116 200 118
rect 194 114 200 116
rect 160 110 166 112
rect 26 85 28 90
rect 36 85 38 90
rect 46 88 48 92
rect 66 85 68 90
rect 76 85 78 90
rect 86 88 88 92
rect 123 88 125 92
rect 133 88 135 92
rect 113 79 115 83
rect 160 108 162 110
rect 164 108 166 110
rect 160 106 166 108
rect 174 110 180 112
rect 174 108 176 110
rect 178 108 180 110
rect 174 106 180 108
rect 178 103 180 106
rect 188 103 190 114
rect 198 110 200 114
rect 231 112 233 125
rect 238 120 240 125
rect 251 120 253 125
rect 237 118 243 120
rect 237 116 239 118
rect 241 116 243 118
rect 237 114 243 116
rect 247 118 253 120
rect 247 116 249 118
rect 251 116 253 118
rect 247 114 253 116
rect 227 110 233 112
rect 227 108 229 110
rect 231 108 233 110
rect 227 106 233 108
rect 231 103 233 106
rect 241 103 243 114
rect 251 110 253 114
rect 271 112 273 125
rect 278 120 280 125
rect 291 120 293 125
rect 277 118 283 120
rect 277 116 279 118
rect 281 116 283 118
rect 277 114 283 116
rect 287 118 293 120
rect 319 119 321 128
rect 326 125 328 128
rect 326 123 330 125
rect 336 124 338 128
rect 346 125 348 128
rect 328 120 330 123
rect 346 123 355 125
rect 403 134 405 138
rect 346 121 351 123
rect 353 121 355 123
rect 287 116 289 118
rect 291 116 293 118
rect 287 114 293 116
rect 267 110 273 112
rect 178 85 180 90
rect 188 85 190 90
rect 198 88 200 92
rect 267 108 269 110
rect 271 108 273 110
rect 267 106 273 108
rect 271 103 273 106
rect 281 103 283 114
rect 291 110 293 114
rect 318 117 324 119
rect 318 115 320 117
rect 322 115 324 117
rect 318 113 324 115
rect 328 118 334 120
rect 328 116 330 118
rect 332 116 334 118
rect 328 114 334 116
rect 346 119 355 121
rect 346 115 348 119
rect 362 115 364 123
rect 318 110 320 113
rect 328 110 330 114
rect 338 113 348 115
rect 354 113 367 115
rect 338 110 340 113
rect 354 110 356 113
rect 365 112 367 113
rect 383 112 385 125
rect 390 120 392 125
rect 403 120 405 125
rect 389 118 395 120
rect 389 116 391 118
rect 393 116 395 118
rect 389 114 395 116
rect 399 118 405 120
rect 399 116 401 118
rect 403 116 405 118
rect 399 114 405 116
rect 365 110 371 112
rect 231 85 233 90
rect 241 85 243 90
rect 251 88 253 92
rect 149 79 151 83
rect 271 85 273 90
rect 281 85 283 90
rect 291 88 293 92
rect 328 88 330 92
rect 338 88 340 92
rect 318 79 320 83
rect 365 108 367 110
rect 369 108 371 110
rect 365 106 371 108
rect 379 110 385 112
rect 379 108 381 110
rect 383 108 385 110
rect 379 106 385 108
rect 383 103 385 106
rect 393 103 395 114
rect 403 110 405 114
rect 383 85 385 90
rect 393 85 395 90
rect 403 88 405 92
rect 354 79 356 83
rect 26 62 28 66
rect 36 64 38 69
rect 46 64 48 69
rect 66 64 68 69
rect 76 64 78 69
rect 155 71 157 75
rect 86 62 88 66
rect 106 62 108 66
rect 116 64 118 69
rect 126 64 128 69
rect 26 40 28 44
rect 36 40 38 51
rect 46 48 48 51
rect 66 48 68 51
rect 46 46 52 48
rect 46 44 48 46
rect 50 44 52 46
rect 46 42 52 44
rect 62 46 68 48
rect 62 44 64 46
rect 66 44 68 46
rect 62 42 68 44
rect 26 38 32 40
rect 26 36 28 38
rect 30 36 32 38
rect 26 34 32 36
rect 36 38 42 40
rect 36 36 38 38
rect 40 36 42 38
rect 36 34 42 36
rect 26 29 28 34
rect 39 29 41 34
rect 46 29 48 42
rect 66 29 68 42
rect 76 40 78 51
rect 86 40 88 44
rect 72 38 78 40
rect 72 36 74 38
rect 76 36 78 38
rect 72 34 78 36
rect 82 38 88 40
rect 82 36 84 38
rect 86 36 88 38
rect 82 34 88 36
rect 73 29 75 34
rect 86 29 88 34
rect 106 40 108 44
rect 116 40 118 51
rect 126 48 128 51
rect 126 46 132 48
rect 126 44 128 46
rect 130 44 132 46
rect 126 42 132 44
rect 140 46 146 48
rect 140 44 142 46
rect 144 44 146 46
rect 191 71 193 75
rect 171 62 173 66
rect 181 62 183 66
rect 231 62 233 66
rect 241 64 243 69
rect 251 64 253 69
rect 271 64 273 69
rect 281 64 283 69
rect 360 71 362 75
rect 291 62 293 66
rect 311 62 313 66
rect 321 64 323 69
rect 331 64 333 69
rect 140 42 146 44
rect 106 38 112 40
rect 106 36 108 38
rect 110 36 112 38
rect 106 34 112 36
rect 116 38 122 40
rect 116 36 118 38
rect 120 36 122 38
rect 116 34 122 36
rect 106 29 108 34
rect 119 29 121 34
rect 126 29 128 42
rect 144 41 146 42
rect 155 41 157 44
rect 171 41 173 44
rect 144 39 157 41
rect 163 39 173 41
rect 181 40 183 44
rect 191 41 193 44
rect 147 31 149 39
rect 163 35 165 39
rect 156 33 165 35
rect 177 38 183 40
rect 177 36 179 38
rect 181 36 183 38
rect 177 34 183 36
rect 187 39 193 41
rect 187 37 189 39
rect 191 37 193 39
rect 187 35 193 37
rect 231 40 233 44
rect 241 40 243 51
rect 251 48 253 51
rect 271 48 273 51
rect 251 46 257 48
rect 251 44 253 46
rect 255 44 257 46
rect 251 42 257 44
rect 267 46 273 48
rect 267 44 269 46
rect 271 44 273 46
rect 267 42 273 44
rect 231 38 237 40
rect 231 36 233 38
rect 235 36 237 38
rect 156 31 158 33
rect 160 31 165 33
rect 26 16 28 20
rect 39 13 41 18
rect 46 13 48 18
rect 66 13 68 18
rect 73 13 75 18
rect 86 16 88 20
rect 106 16 108 20
rect 156 29 165 31
rect 181 31 183 34
rect 163 26 165 29
rect 173 26 175 30
rect 181 29 185 31
rect 183 26 185 29
rect 190 26 192 35
rect 231 34 237 36
rect 241 38 247 40
rect 241 36 243 38
rect 245 36 247 38
rect 241 34 247 36
rect 231 29 233 34
rect 244 29 246 34
rect 251 29 253 42
rect 271 29 273 42
rect 281 40 283 51
rect 291 40 293 44
rect 277 38 283 40
rect 277 36 279 38
rect 281 36 283 38
rect 277 34 283 36
rect 287 38 293 40
rect 287 36 289 38
rect 291 36 293 38
rect 287 34 293 36
rect 278 29 280 34
rect 291 29 293 34
rect 311 40 313 44
rect 321 40 323 51
rect 331 48 333 51
rect 331 46 337 48
rect 331 44 333 46
rect 335 44 337 46
rect 331 42 337 44
rect 345 46 351 48
rect 345 44 347 46
rect 349 44 351 46
rect 396 71 398 75
rect 376 62 378 66
rect 386 62 388 66
rect 345 42 351 44
rect 311 38 317 40
rect 311 36 313 38
rect 315 36 317 38
rect 311 34 317 36
rect 321 38 327 40
rect 321 36 323 38
rect 325 36 327 38
rect 321 34 327 36
rect 311 29 313 34
rect 324 29 326 34
rect 331 29 333 42
rect 349 41 351 42
rect 360 41 362 44
rect 376 41 378 44
rect 349 39 362 41
rect 368 39 378 41
rect 386 40 388 44
rect 396 41 398 44
rect 352 31 354 39
rect 368 35 370 39
rect 361 33 370 35
rect 382 38 388 40
rect 382 36 384 38
rect 386 36 388 38
rect 382 34 388 36
rect 392 39 398 41
rect 392 37 394 39
rect 396 37 398 39
rect 392 35 398 37
rect 361 31 363 33
rect 365 31 370 33
rect 147 19 149 22
rect 119 13 121 18
rect 126 13 128 18
rect 147 17 152 19
rect 150 9 152 17
rect 163 13 165 17
rect 173 9 175 17
rect 231 16 233 20
rect 183 9 185 14
rect 190 9 192 14
rect 150 7 175 9
rect 244 13 246 18
rect 251 13 253 18
rect 271 13 273 18
rect 278 13 280 18
rect 291 16 293 20
rect 311 16 313 20
rect 361 29 370 31
rect 386 31 388 34
rect 368 26 370 29
rect 378 26 380 30
rect 386 29 390 31
rect 388 26 390 29
rect 395 26 397 35
rect 352 19 354 22
rect 324 13 326 18
rect 331 13 333 18
rect 352 17 357 19
rect 355 9 357 17
rect 368 13 370 17
rect 378 9 380 17
rect 388 9 390 14
rect 395 9 397 14
rect 355 7 380 9
rect -240 -12 -238 -7
rect -230 -15 -228 -10
rect -220 -15 -218 -10
rect -200 -10 -198 -6
rect -187 -8 -185 -3
rect -180 -8 -178 -3
rect -156 1 -131 3
rect -156 -7 -154 1
rect -143 -7 -141 -3
rect -133 -7 -131 1
rect -123 -4 -121 1
rect -116 -4 -114 1
rect -159 -9 -154 -7
rect -159 -12 -157 -9
rect -240 -24 -238 -21
rect -230 -24 -228 -21
rect -240 -26 -234 -24
rect -240 -28 -238 -26
rect -236 -28 -234 -26
rect -240 -30 -234 -28
rect -230 -26 -224 -24
rect -230 -28 -228 -26
rect -226 -28 -224 -26
rect -230 -30 -224 -28
rect -240 -33 -238 -30
rect -227 -40 -225 -30
rect -220 -31 -218 -21
rect -200 -24 -198 -19
rect -187 -24 -185 -19
rect -200 -26 -194 -24
rect -200 -28 -198 -26
rect -196 -28 -194 -26
rect -200 -30 -194 -28
rect -190 -26 -184 -24
rect -190 -28 -188 -26
rect -186 -28 -184 -26
rect -190 -30 -184 -28
rect -220 -33 -214 -31
rect -220 -35 -218 -33
rect -216 -35 -214 -33
rect -200 -34 -198 -30
rect -220 -37 -214 -35
rect -220 -40 -218 -37
rect -240 -56 -238 -51
rect -190 -41 -188 -30
rect -180 -32 -178 -19
rect -95 -10 -93 -6
rect -82 -8 -80 -3
rect -75 -8 -73 -3
rect -51 1 -26 3
rect -51 -7 -49 1
rect -38 -7 -36 -3
rect -28 -7 -26 1
rect -18 -4 -16 1
rect -11 -4 -9 1
rect -143 -19 -141 -16
rect -150 -21 -141 -19
rect -133 -20 -131 -16
rect -123 -19 -121 -16
rect -159 -29 -157 -21
rect -150 -23 -148 -21
rect -146 -23 -141 -21
rect -150 -25 -141 -23
rect -125 -21 -121 -19
rect -125 -24 -123 -21
rect -143 -29 -141 -25
rect -129 -26 -123 -24
rect -116 -25 -114 -16
rect -54 -9 -49 -7
rect -54 -12 -52 -9
rect -95 -24 -93 -19
rect -82 -24 -80 -19
rect -129 -28 -127 -26
rect -125 -28 -123 -26
rect -162 -31 -149 -29
rect -143 -31 -133 -29
rect -129 -30 -123 -28
rect -162 -32 -160 -31
rect -180 -34 -174 -32
rect -180 -36 -178 -34
rect -176 -36 -174 -34
rect -180 -38 -174 -36
rect -166 -34 -160 -32
rect -151 -34 -149 -31
rect -135 -34 -133 -31
rect -125 -34 -123 -30
rect -119 -27 -113 -25
rect -119 -29 -117 -27
rect -115 -29 -113 -27
rect -119 -31 -113 -29
rect -115 -34 -113 -31
rect -95 -26 -89 -24
rect -95 -28 -93 -26
rect -91 -28 -89 -26
rect -95 -30 -89 -28
rect -85 -26 -79 -24
rect -85 -28 -83 -26
rect -81 -28 -79 -26
rect -85 -30 -79 -28
rect -95 -34 -93 -30
rect -166 -36 -164 -34
rect -162 -36 -160 -34
rect -166 -38 -160 -36
rect -180 -41 -178 -38
rect -200 -56 -198 -52
rect -190 -59 -188 -54
rect -180 -59 -178 -54
rect -227 -65 -225 -61
rect -220 -65 -218 -61
rect -135 -56 -133 -52
rect -125 -56 -123 -52
rect -151 -65 -149 -61
rect -85 -41 -83 -30
rect -75 -32 -73 -19
rect 10 -12 12 -7
rect -38 -19 -36 -16
rect -45 -21 -36 -19
rect -28 -20 -26 -16
rect -18 -19 -16 -16
rect -54 -29 -52 -21
rect -45 -23 -43 -21
rect -41 -23 -36 -21
rect -45 -25 -36 -23
rect -20 -21 -16 -19
rect -20 -24 -18 -21
rect -38 -29 -36 -25
rect -24 -26 -18 -24
rect -11 -25 -9 -16
rect 20 -15 22 -10
rect 30 -15 32 -10
rect 50 -10 52 -6
rect 63 -8 65 -3
rect 70 -8 72 -3
rect 94 1 119 3
rect 94 -7 96 1
rect 107 -7 109 -3
rect 117 -7 119 1
rect 127 -4 129 1
rect 134 -4 136 1
rect 91 -9 96 -7
rect 91 -12 93 -9
rect 10 -24 12 -21
rect 20 -24 22 -21
rect -24 -28 -22 -26
rect -20 -28 -18 -26
rect -57 -31 -44 -29
rect -38 -31 -28 -29
rect -24 -30 -18 -28
rect -57 -32 -55 -31
rect -75 -34 -69 -32
rect -75 -36 -73 -34
rect -71 -36 -69 -34
rect -75 -38 -69 -36
rect -61 -34 -55 -32
rect -46 -34 -44 -31
rect -30 -34 -28 -31
rect -20 -34 -18 -30
rect -14 -27 -8 -25
rect -14 -29 -12 -27
rect -10 -29 -8 -27
rect -14 -31 -8 -29
rect -10 -34 -8 -31
rect 10 -26 16 -24
rect 10 -28 12 -26
rect 14 -28 16 -26
rect 10 -30 16 -28
rect 20 -26 26 -24
rect 20 -28 22 -26
rect 24 -28 26 -26
rect 20 -30 26 -28
rect 10 -33 12 -30
rect -61 -36 -59 -34
rect -57 -36 -55 -34
rect -61 -38 -55 -36
rect -75 -41 -73 -38
rect -95 -56 -93 -52
rect -85 -59 -83 -54
rect -75 -59 -73 -54
rect -115 -65 -113 -61
rect -30 -56 -28 -52
rect -20 -56 -18 -52
rect -46 -65 -44 -61
rect 23 -40 25 -30
rect 30 -31 32 -21
rect 50 -24 52 -19
rect 63 -24 65 -19
rect 50 -26 56 -24
rect 50 -28 52 -26
rect 54 -28 56 -26
rect 50 -30 56 -28
rect 60 -26 66 -24
rect 60 -28 62 -26
rect 64 -28 66 -26
rect 60 -30 66 -28
rect 30 -33 36 -31
rect 30 -35 32 -33
rect 34 -35 36 -33
rect 50 -34 52 -30
rect 30 -37 36 -35
rect 30 -40 32 -37
rect 10 -56 12 -51
rect -10 -65 -8 -61
rect 60 -41 62 -30
rect 70 -32 72 -19
rect 155 -10 157 -6
rect 168 -8 170 -3
rect 175 -8 177 -3
rect 199 1 224 3
rect 199 -7 201 1
rect 212 -7 214 -3
rect 222 -7 224 1
rect 232 -4 234 1
rect 239 -4 241 1
rect 107 -19 109 -16
rect 100 -21 109 -19
rect 117 -20 119 -16
rect 127 -19 129 -16
rect 91 -29 93 -21
rect 100 -23 102 -21
rect 104 -23 109 -21
rect 100 -25 109 -23
rect 125 -21 129 -19
rect 125 -24 127 -21
rect 107 -29 109 -25
rect 121 -26 127 -24
rect 134 -25 136 -16
rect 196 -9 201 -7
rect 196 -12 198 -9
rect 155 -24 157 -19
rect 168 -24 170 -19
rect 121 -28 123 -26
rect 125 -28 127 -26
rect 88 -31 101 -29
rect 107 -31 117 -29
rect 121 -30 127 -28
rect 88 -32 90 -31
rect 70 -34 76 -32
rect 70 -36 72 -34
rect 74 -36 76 -34
rect 70 -38 76 -36
rect 84 -34 90 -32
rect 99 -34 101 -31
rect 115 -34 117 -31
rect 125 -34 127 -30
rect 131 -27 137 -25
rect 131 -29 133 -27
rect 135 -29 137 -27
rect 131 -31 137 -29
rect 135 -34 137 -31
rect 155 -26 161 -24
rect 155 -28 157 -26
rect 159 -28 161 -26
rect 155 -30 161 -28
rect 165 -26 171 -24
rect 165 -28 167 -26
rect 169 -28 171 -26
rect 165 -30 171 -28
rect 155 -34 157 -30
rect 84 -36 86 -34
rect 88 -36 90 -34
rect 84 -38 90 -36
rect 70 -41 72 -38
rect 50 -56 52 -52
rect 60 -59 62 -54
rect 70 -59 72 -54
rect 23 -65 25 -61
rect 30 -65 32 -61
rect 115 -56 117 -52
rect 125 -56 127 -52
rect 99 -65 101 -61
rect 165 -41 167 -30
rect 175 -32 177 -19
rect 260 -12 262 -7
rect 212 -19 214 -16
rect 205 -21 214 -19
rect 222 -20 224 -16
rect 232 -19 234 -16
rect 196 -29 198 -21
rect 205 -23 207 -21
rect 209 -23 214 -21
rect 205 -25 214 -23
rect 230 -21 234 -19
rect 230 -24 232 -21
rect 212 -29 214 -25
rect 226 -26 232 -24
rect 239 -25 241 -16
rect 270 -15 272 -10
rect 280 -15 282 -10
rect 300 -10 302 -6
rect 313 -8 315 -3
rect 320 -8 322 -3
rect 344 1 369 3
rect 344 -7 346 1
rect 357 -7 359 -3
rect 367 -7 369 1
rect 377 -4 379 1
rect 384 -4 386 1
rect 341 -9 346 -7
rect 341 -12 343 -9
rect 260 -24 262 -21
rect 270 -24 272 -21
rect 226 -28 228 -26
rect 230 -28 232 -26
rect 193 -31 206 -29
rect 212 -31 222 -29
rect 226 -30 232 -28
rect 193 -32 195 -31
rect 175 -34 181 -32
rect 175 -36 177 -34
rect 179 -36 181 -34
rect 175 -38 181 -36
rect 189 -34 195 -32
rect 204 -34 206 -31
rect 220 -34 222 -31
rect 230 -34 232 -30
rect 236 -27 242 -25
rect 236 -29 238 -27
rect 240 -29 242 -27
rect 236 -31 242 -29
rect 240 -34 242 -31
rect 260 -26 266 -24
rect 260 -28 262 -26
rect 264 -28 266 -26
rect 260 -30 266 -28
rect 270 -26 276 -24
rect 270 -28 272 -26
rect 274 -28 276 -26
rect 270 -30 276 -28
rect 260 -33 262 -30
rect 189 -36 191 -34
rect 193 -36 195 -34
rect 189 -38 195 -36
rect 175 -41 177 -38
rect 155 -56 157 -52
rect 165 -59 167 -54
rect 175 -59 177 -54
rect 135 -65 137 -61
rect 220 -56 222 -52
rect 230 -56 232 -52
rect 204 -65 206 -61
rect 273 -40 275 -30
rect 280 -31 282 -21
rect 300 -24 302 -19
rect 313 -24 315 -19
rect 300 -26 306 -24
rect 300 -28 302 -26
rect 304 -28 306 -26
rect 300 -30 306 -28
rect 310 -26 316 -24
rect 310 -28 312 -26
rect 314 -28 316 -26
rect 310 -30 316 -28
rect 280 -33 286 -31
rect 280 -35 282 -33
rect 284 -35 286 -33
rect 300 -34 302 -30
rect 280 -37 286 -35
rect 280 -40 282 -37
rect 260 -56 262 -51
rect 240 -65 242 -61
rect 310 -41 312 -30
rect 320 -32 322 -19
rect 405 -10 407 -6
rect 418 -8 420 -3
rect 425 -8 427 -3
rect 449 1 474 3
rect 449 -7 451 1
rect 462 -7 464 -3
rect 472 -7 474 1
rect 482 -4 484 1
rect 489 -4 491 1
rect 357 -19 359 -16
rect 350 -21 359 -19
rect 367 -20 369 -16
rect 377 -19 379 -16
rect 341 -29 343 -21
rect 350 -23 352 -21
rect 354 -23 359 -21
rect 350 -25 359 -23
rect 375 -21 379 -19
rect 375 -24 377 -21
rect 357 -29 359 -25
rect 371 -26 377 -24
rect 384 -25 386 -16
rect 446 -9 451 -7
rect 446 -12 448 -9
rect 405 -24 407 -19
rect 418 -24 420 -19
rect 371 -28 373 -26
rect 375 -28 377 -26
rect 338 -31 351 -29
rect 357 -31 367 -29
rect 371 -30 377 -28
rect 338 -32 340 -31
rect 320 -34 326 -32
rect 320 -36 322 -34
rect 324 -36 326 -34
rect 320 -38 326 -36
rect 334 -34 340 -32
rect 349 -34 351 -31
rect 365 -34 367 -31
rect 375 -34 377 -30
rect 381 -27 387 -25
rect 381 -29 383 -27
rect 385 -29 387 -27
rect 381 -31 387 -29
rect 385 -34 387 -31
rect 405 -26 411 -24
rect 405 -28 407 -26
rect 409 -28 411 -26
rect 405 -30 411 -28
rect 415 -26 421 -24
rect 415 -28 417 -26
rect 419 -28 421 -26
rect 415 -30 421 -28
rect 405 -34 407 -30
rect 334 -36 336 -34
rect 338 -36 340 -34
rect 334 -38 340 -36
rect 320 -41 322 -38
rect 300 -56 302 -52
rect 310 -59 312 -54
rect 320 -59 322 -54
rect 273 -65 275 -61
rect 280 -65 282 -61
rect 365 -56 367 -52
rect 375 -56 377 -52
rect 349 -65 351 -61
rect 415 -41 417 -30
rect 425 -32 427 -19
rect 510 -12 512 -7
rect 462 -19 464 -16
rect 455 -21 464 -19
rect 472 -20 474 -16
rect 482 -19 484 -16
rect 446 -29 448 -21
rect 455 -23 457 -21
rect 459 -23 464 -21
rect 455 -25 464 -23
rect 480 -21 484 -19
rect 480 -24 482 -21
rect 462 -29 464 -25
rect 476 -26 482 -24
rect 489 -25 491 -16
rect 520 -15 522 -10
rect 530 -15 532 -10
rect 550 -10 552 -6
rect 563 -8 565 -3
rect 570 -8 572 -3
rect 594 1 619 3
rect 594 -7 596 1
rect 607 -7 609 -3
rect 617 -7 619 1
rect 627 -4 629 1
rect 634 -4 636 1
rect 591 -9 596 -7
rect 591 -12 593 -9
rect 510 -24 512 -21
rect 520 -24 522 -21
rect 476 -28 478 -26
rect 480 -28 482 -26
rect 443 -31 456 -29
rect 462 -31 472 -29
rect 476 -30 482 -28
rect 443 -32 445 -31
rect 425 -34 431 -32
rect 425 -36 427 -34
rect 429 -36 431 -34
rect 425 -38 431 -36
rect 439 -34 445 -32
rect 454 -34 456 -31
rect 470 -34 472 -31
rect 480 -34 482 -30
rect 486 -27 492 -25
rect 486 -29 488 -27
rect 490 -29 492 -27
rect 486 -31 492 -29
rect 490 -34 492 -31
rect 510 -26 516 -24
rect 510 -28 512 -26
rect 514 -28 516 -26
rect 510 -30 516 -28
rect 520 -26 526 -24
rect 520 -28 522 -26
rect 524 -28 526 -26
rect 520 -30 526 -28
rect 510 -33 512 -30
rect 439 -36 441 -34
rect 443 -36 445 -34
rect 439 -38 445 -36
rect 425 -41 427 -38
rect 405 -56 407 -52
rect 415 -59 417 -54
rect 425 -59 427 -54
rect 385 -65 387 -61
rect 470 -56 472 -52
rect 480 -56 482 -52
rect 454 -65 456 -61
rect 523 -40 525 -30
rect 530 -31 532 -21
rect 550 -24 552 -19
rect 563 -24 565 -19
rect 550 -26 556 -24
rect 550 -28 552 -26
rect 554 -28 556 -26
rect 550 -30 556 -28
rect 560 -26 566 -24
rect 560 -28 562 -26
rect 564 -28 566 -26
rect 560 -30 566 -28
rect 530 -33 536 -31
rect 530 -35 532 -33
rect 534 -35 536 -33
rect 550 -34 552 -30
rect 530 -37 536 -35
rect 530 -40 532 -37
rect 510 -56 512 -51
rect 490 -65 492 -61
rect 560 -41 562 -30
rect 570 -32 572 -19
rect 655 -10 657 -6
rect 668 -8 670 -3
rect 675 -8 677 -3
rect 699 1 724 3
rect 699 -7 701 1
rect 712 -7 714 -3
rect 722 -7 724 1
rect 732 -4 734 1
rect 739 -4 741 1
rect 607 -19 609 -16
rect 600 -21 609 -19
rect 617 -20 619 -16
rect 627 -19 629 -16
rect 591 -29 593 -21
rect 600 -23 602 -21
rect 604 -23 609 -21
rect 600 -25 609 -23
rect 625 -21 629 -19
rect 625 -24 627 -21
rect 607 -29 609 -25
rect 621 -26 627 -24
rect 634 -25 636 -16
rect 696 -9 701 -7
rect 696 -12 698 -9
rect 655 -24 657 -19
rect 668 -24 670 -19
rect 621 -28 623 -26
rect 625 -28 627 -26
rect 588 -31 601 -29
rect 607 -31 617 -29
rect 621 -30 627 -28
rect 588 -32 590 -31
rect 570 -34 576 -32
rect 570 -36 572 -34
rect 574 -36 576 -34
rect 570 -38 576 -36
rect 584 -34 590 -32
rect 599 -34 601 -31
rect 615 -34 617 -31
rect 625 -34 627 -30
rect 631 -27 637 -25
rect 631 -29 633 -27
rect 635 -29 637 -27
rect 631 -31 637 -29
rect 635 -34 637 -31
rect 655 -26 661 -24
rect 655 -28 657 -26
rect 659 -28 661 -26
rect 655 -30 661 -28
rect 665 -26 671 -24
rect 665 -28 667 -26
rect 669 -28 671 -26
rect 665 -30 671 -28
rect 655 -34 657 -30
rect 584 -36 586 -34
rect 588 -36 590 -34
rect 584 -38 590 -36
rect 570 -41 572 -38
rect 550 -56 552 -52
rect 560 -59 562 -54
rect 570 -59 572 -54
rect 523 -65 525 -61
rect 530 -65 532 -61
rect 615 -56 617 -52
rect 625 -56 627 -52
rect 599 -65 601 -61
rect 665 -41 667 -30
rect 675 -32 677 -19
rect 712 -19 714 -16
rect 705 -21 714 -19
rect 722 -20 724 -16
rect 732 -19 734 -16
rect 696 -29 698 -21
rect 705 -23 707 -21
rect 709 -23 714 -21
rect 705 -25 714 -23
rect 730 -21 734 -19
rect 730 -24 732 -21
rect 712 -29 714 -25
rect 726 -26 732 -24
rect 739 -25 741 -16
rect 726 -28 728 -26
rect 730 -28 732 -26
rect 693 -31 706 -29
rect 712 -31 722 -29
rect 726 -30 732 -28
rect 693 -32 695 -31
rect 675 -34 681 -32
rect 675 -36 677 -34
rect 679 -36 681 -34
rect 675 -38 681 -36
rect 689 -34 695 -32
rect 704 -34 706 -31
rect 720 -34 722 -31
rect 730 -34 732 -30
rect 736 -27 742 -25
rect 736 -29 738 -27
rect 740 -29 742 -27
rect 736 -31 742 -29
rect 740 -34 742 -31
rect 689 -36 691 -34
rect 693 -36 695 -34
rect 689 -38 695 -36
rect 675 -41 677 -38
rect 655 -56 657 -52
rect 665 -59 667 -54
rect 675 -59 677 -54
rect 635 -65 637 -61
rect 720 -56 722 -52
rect 730 -56 732 -52
rect 704 -65 706 -61
rect 740 -65 742 -61
<< ndif >>
rect 37 144 44 146
rect 37 142 40 144
rect 42 142 44 144
rect 37 136 44 142
rect 77 144 84 146
rect 77 142 80 144
rect 82 142 84 144
rect 19 134 26 136
rect 19 132 21 134
rect 23 132 26 134
rect 19 130 26 132
rect 21 125 26 130
rect 28 125 33 136
rect 35 134 44 136
rect 77 136 84 142
rect 106 144 112 146
rect 106 142 108 144
rect 110 142 112 144
rect 106 140 112 142
rect 59 134 66 136
rect 35 125 46 134
rect 48 132 55 134
rect 48 130 51 132
rect 53 130 55 132
rect 59 132 61 134
rect 63 132 66 134
rect 59 130 66 132
rect 48 128 55 130
rect 48 125 53 128
rect 61 125 66 130
rect 68 125 73 136
rect 75 134 84 136
rect 75 125 86 134
rect 88 132 95 134
rect 88 130 91 132
rect 93 130 95 132
rect 88 128 95 130
rect 106 128 114 140
rect 116 128 121 140
rect 123 137 128 140
rect 189 144 196 146
rect 189 142 192 144
rect 194 142 196 144
rect 123 134 131 137
rect 123 132 126 134
rect 128 132 131 134
rect 123 128 131 132
rect 133 132 141 137
rect 133 130 136 132
rect 138 130 141 132
rect 133 128 141 130
rect 143 135 152 137
rect 189 136 196 142
rect 242 144 249 146
rect 242 142 245 144
rect 247 142 249 144
rect 143 133 148 135
rect 150 133 152 135
rect 143 132 152 133
rect 171 134 178 136
rect 171 132 173 134
rect 175 132 178 134
rect 143 128 157 132
rect 88 125 93 128
rect 152 123 157 128
rect 159 129 164 132
rect 171 130 178 132
rect 159 127 166 129
rect 159 125 162 127
rect 164 125 166 127
rect 173 125 178 130
rect 180 125 185 136
rect 187 134 196 136
rect 242 136 249 142
rect 282 144 289 146
rect 282 142 285 144
rect 287 142 289 144
rect 224 134 231 136
rect 187 125 198 134
rect 200 132 207 134
rect 200 130 203 132
rect 205 130 207 132
rect 224 132 226 134
rect 228 132 231 134
rect 224 130 231 132
rect 200 128 207 130
rect 200 125 205 128
rect 226 125 231 130
rect 233 125 238 136
rect 240 134 249 136
rect 282 136 289 142
rect 311 144 317 146
rect 311 142 313 144
rect 315 142 317 144
rect 311 140 317 142
rect 264 134 271 136
rect 240 125 251 134
rect 253 132 260 134
rect 253 130 256 132
rect 258 130 260 132
rect 264 132 266 134
rect 268 132 271 134
rect 264 130 271 132
rect 253 128 260 130
rect 253 125 258 128
rect 266 125 271 130
rect 273 125 278 136
rect 280 134 289 136
rect 280 125 291 134
rect 293 132 300 134
rect 293 130 296 132
rect 298 130 300 132
rect 293 128 300 130
rect 311 128 319 140
rect 321 128 326 140
rect 328 137 333 140
rect 394 144 401 146
rect 394 142 397 144
rect 399 142 401 144
rect 328 134 336 137
rect 328 132 331 134
rect 333 132 336 134
rect 328 128 336 132
rect 338 132 346 137
rect 338 130 341 132
rect 343 130 346 132
rect 338 128 346 130
rect 348 135 357 137
rect 394 136 401 142
rect 348 133 353 135
rect 355 133 357 135
rect 348 132 357 133
rect 376 134 383 136
rect 376 132 378 134
rect 380 132 383 134
rect 348 128 362 132
rect 293 125 298 128
rect 159 123 166 125
rect 357 123 362 128
rect 364 129 369 132
rect 376 130 383 132
rect 364 127 371 129
rect 364 125 367 127
rect 369 125 371 127
rect 378 125 383 130
rect 385 125 390 136
rect 392 134 401 136
rect 392 125 403 134
rect 405 132 412 134
rect 405 130 408 132
rect 410 130 412 132
rect 405 128 412 130
rect 405 125 410 128
rect 364 123 371 125
rect 140 29 147 31
rect 21 26 26 29
rect 19 24 26 26
rect 19 22 21 24
rect 23 22 26 24
rect 19 20 26 22
rect 28 20 39 29
rect 30 18 39 20
rect 41 18 46 29
rect 48 24 53 29
rect 61 24 66 29
rect 48 22 55 24
rect 48 20 51 22
rect 53 20 55 22
rect 48 18 55 20
rect 59 22 66 24
rect 59 20 61 22
rect 63 20 66 22
rect 59 18 66 20
rect 68 18 73 29
rect 75 20 86 29
rect 88 26 93 29
rect 101 26 106 29
rect 88 24 95 26
rect 88 22 91 24
rect 93 22 95 24
rect 88 20 95 22
rect 99 24 106 26
rect 99 22 101 24
rect 103 22 106 24
rect 99 20 106 22
rect 108 20 119 29
rect 75 18 84 20
rect 30 12 37 18
rect 30 10 32 12
rect 34 10 37 12
rect 30 8 37 10
rect 77 12 84 18
rect 110 18 119 20
rect 121 18 126 29
rect 128 24 133 29
rect 140 27 142 29
rect 144 27 147 29
rect 140 25 147 27
rect 128 22 135 24
rect 142 22 147 25
rect 149 26 154 31
rect 345 29 352 31
rect 226 26 231 29
rect 149 22 163 26
rect 128 20 131 22
rect 133 20 135 22
rect 128 18 135 20
rect 154 21 163 22
rect 154 19 156 21
rect 158 19 163 21
rect 77 10 80 12
rect 82 10 84 12
rect 77 8 84 10
rect 110 12 117 18
rect 154 17 163 19
rect 165 24 173 26
rect 165 22 168 24
rect 170 22 173 24
rect 165 17 173 22
rect 175 22 183 26
rect 175 20 178 22
rect 180 20 183 22
rect 175 17 183 20
rect 110 10 112 12
rect 114 10 117 12
rect 110 8 117 10
rect 178 14 183 17
rect 185 14 190 26
rect 192 14 200 26
rect 224 24 231 26
rect 224 22 226 24
rect 228 22 231 24
rect 224 20 231 22
rect 233 20 244 29
rect 235 18 244 20
rect 246 18 251 29
rect 253 24 258 29
rect 266 24 271 29
rect 253 22 260 24
rect 253 20 256 22
rect 258 20 260 22
rect 253 18 260 20
rect 264 22 271 24
rect 264 20 266 22
rect 268 20 271 22
rect 264 18 271 20
rect 273 18 278 29
rect 280 20 291 29
rect 293 26 298 29
rect 306 26 311 29
rect 293 24 300 26
rect 293 22 296 24
rect 298 22 300 24
rect 293 20 300 22
rect 304 24 311 26
rect 304 22 306 24
rect 308 22 311 24
rect 304 20 311 22
rect 313 20 324 29
rect 280 18 289 20
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
rect 235 12 242 18
rect 235 10 237 12
rect 239 10 242 12
rect 235 8 242 10
rect 282 12 289 18
rect 315 18 324 20
rect 326 18 331 29
rect 333 24 338 29
rect 345 27 347 29
rect 349 27 352 29
rect 345 25 352 27
rect 333 22 340 24
rect 347 22 352 25
rect 354 26 359 31
rect 354 22 368 26
rect 333 20 336 22
rect 338 20 340 22
rect 333 18 340 20
rect 359 21 368 22
rect 359 19 361 21
rect 363 19 368 21
rect 282 10 285 12
rect 287 10 289 12
rect 282 8 289 10
rect 315 12 322 18
rect 359 17 368 19
rect 370 24 378 26
rect 370 22 373 24
rect 375 22 378 24
rect 370 17 378 22
rect 380 22 388 26
rect 380 20 383 22
rect 385 20 388 22
rect 380 17 388 20
rect 315 10 317 12
rect 319 10 322 12
rect 315 8 322 10
rect 383 14 388 17
rect 390 14 395 26
rect 397 14 405 26
rect 399 12 405 14
rect 399 10 401 12
rect 403 10 405 12
rect 399 8 405 10
rect -236 -4 -230 -2
rect -236 -6 -234 -4
rect -232 -6 -230 -4
rect -236 -8 -230 -6
rect -217 -4 -211 -2
rect -196 0 -189 2
rect -196 -2 -194 0
rect -192 -2 -189 0
rect -217 -6 -215 -4
rect -213 -6 -211 -4
rect -217 -8 -211 -6
rect -236 -12 -232 -8
rect -245 -15 -240 -12
rect -247 -17 -240 -15
rect -247 -19 -245 -17
rect -243 -19 -240 -17
rect -247 -21 -240 -19
rect -238 -15 -232 -12
rect -216 -15 -211 -8
rect -196 -8 -189 -2
rect -112 0 -106 2
rect -112 -2 -110 0
rect -108 -2 -106 0
rect -112 -4 -106 -2
rect -91 0 -84 2
rect -91 -2 -89 0
rect -87 -2 -84 0
rect -128 -7 -123 -4
rect -196 -10 -187 -8
rect -238 -21 -230 -15
rect -228 -17 -220 -15
rect -228 -19 -225 -17
rect -223 -19 -220 -17
rect -228 -21 -220 -19
rect -218 -21 -211 -15
rect -207 -12 -200 -10
rect -207 -14 -205 -12
rect -203 -14 -200 -12
rect -207 -16 -200 -14
rect -205 -19 -200 -16
rect -198 -19 -187 -10
rect -185 -19 -180 -8
rect -178 -10 -171 -8
rect -178 -12 -175 -10
rect -173 -12 -171 -10
rect -152 -9 -143 -7
rect -152 -11 -150 -9
rect -148 -11 -143 -9
rect -152 -12 -143 -11
rect -178 -14 -171 -12
rect -178 -19 -173 -14
rect -164 -15 -159 -12
rect -166 -17 -159 -15
rect -166 -19 -164 -17
rect -162 -19 -159 -17
rect -166 -21 -159 -19
rect -157 -16 -143 -12
rect -141 -12 -133 -7
rect -141 -14 -138 -12
rect -136 -14 -133 -12
rect -141 -16 -133 -14
rect -131 -10 -123 -7
rect -131 -12 -128 -10
rect -126 -12 -123 -10
rect -131 -16 -123 -12
rect -121 -16 -116 -4
rect -114 -16 -106 -4
rect -91 -8 -84 -2
rect -7 0 -1 2
rect -7 -2 -5 0
rect -3 -2 -1 0
rect -7 -4 -1 -2
rect 14 -4 20 -2
rect -23 -7 -18 -4
rect -91 -10 -82 -8
rect -102 -12 -95 -10
rect -102 -14 -100 -12
rect -98 -14 -95 -12
rect -102 -16 -95 -14
rect -157 -21 -152 -16
rect -100 -19 -95 -16
rect -93 -19 -82 -10
rect -80 -19 -75 -8
rect -73 -10 -66 -8
rect -73 -12 -70 -10
rect -68 -12 -66 -10
rect -47 -9 -38 -7
rect -47 -11 -45 -9
rect -43 -11 -38 -9
rect -47 -12 -38 -11
rect -73 -14 -66 -12
rect -73 -19 -68 -14
rect -59 -15 -54 -12
rect -61 -17 -54 -15
rect -61 -19 -59 -17
rect -57 -19 -54 -17
rect -61 -21 -54 -19
rect -52 -16 -38 -12
rect -36 -12 -28 -7
rect -36 -14 -33 -12
rect -31 -14 -28 -12
rect -36 -16 -28 -14
rect -26 -10 -18 -7
rect -26 -12 -23 -10
rect -21 -12 -18 -10
rect -26 -16 -18 -12
rect -16 -16 -11 -4
rect -9 -16 -1 -4
rect 14 -6 16 -4
rect 18 -6 20 -4
rect 14 -8 20 -6
rect 33 -4 39 -2
rect 54 0 61 2
rect 54 -2 56 0
rect 58 -2 61 0
rect 33 -6 35 -4
rect 37 -6 39 -4
rect 33 -8 39 -6
rect 14 -12 18 -8
rect 5 -15 10 -12
rect -52 -21 -47 -16
rect 3 -17 10 -15
rect 3 -19 5 -17
rect 7 -19 10 -17
rect 3 -21 10 -19
rect 12 -15 18 -12
rect 34 -15 39 -8
rect 54 -8 61 -2
rect 138 0 144 2
rect 138 -2 140 0
rect 142 -2 144 0
rect 138 -4 144 -2
rect 159 0 166 2
rect 159 -2 161 0
rect 163 -2 166 0
rect 122 -7 127 -4
rect 54 -10 63 -8
rect 12 -21 20 -15
rect 22 -17 30 -15
rect 22 -19 25 -17
rect 27 -19 30 -17
rect 22 -21 30 -19
rect 32 -21 39 -15
rect 43 -12 50 -10
rect 43 -14 45 -12
rect 47 -14 50 -12
rect 43 -16 50 -14
rect 45 -19 50 -16
rect 52 -19 63 -10
rect 65 -19 70 -8
rect 72 -10 79 -8
rect 72 -12 75 -10
rect 77 -12 79 -10
rect 98 -9 107 -7
rect 98 -11 100 -9
rect 102 -11 107 -9
rect 98 -12 107 -11
rect 72 -14 79 -12
rect 72 -19 77 -14
rect 86 -15 91 -12
rect 84 -17 91 -15
rect 84 -19 86 -17
rect 88 -19 91 -17
rect 84 -21 91 -19
rect 93 -16 107 -12
rect 109 -12 117 -7
rect 109 -14 112 -12
rect 114 -14 117 -12
rect 109 -16 117 -14
rect 119 -10 127 -7
rect 119 -12 122 -10
rect 124 -12 127 -10
rect 119 -16 127 -12
rect 129 -16 134 -4
rect 136 -16 144 -4
rect 159 -8 166 -2
rect 243 0 249 2
rect 243 -2 245 0
rect 247 -2 249 0
rect 243 -4 249 -2
rect 264 -4 270 -2
rect 227 -7 232 -4
rect 159 -10 168 -8
rect 148 -12 155 -10
rect 148 -14 150 -12
rect 152 -14 155 -12
rect 148 -16 155 -14
rect 93 -21 98 -16
rect 150 -19 155 -16
rect 157 -19 168 -10
rect 170 -19 175 -8
rect 177 -10 184 -8
rect 177 -12 180 -10
rect 182 -12 184 -10
rect 203 -9 212 -7
rect 203 -11 205 -9
rect 207 -11 212 -9
rect 203 -12 212 -11
rect 177 -14 184 -12
rect 177 -19 182 -14
rect 191 -15 196 -12
rect 189 -17 196 -15
rect 189 -19 191 -17
rect 193 -19 196 -17
rect 189 -21 196 -19
rect 198 -16 212 -12
rect 214 -12 222 -7
rect 214 -14 217 -12
rect 219 -14 222 -12
rect 214 -16 222 -14
rect 224 -10 232 -7
rect 224 -12 227 -10
rect 229 -12 232 -10
rect 224 -16 232 -12
rect 234 -16 239 -4
rect 241 -16 249 -4
rect 264 -6 266 -4
rect 268 -6 270 -4
rect 264 -8 270 -6
rect 283 -4 289 -2
rect 304 0 311 2
rect 304 -2 306 0
rect 308 -2 311 0
rect 283 -6 285 -4
rect 287 -6 289 -4
rect 283 -8 289 -6
rect 264 -12 268 -8
rect 255 -15 260 -12
rect 198 -21 203 -16
rect 253 -17 260 -15
rect 253 -19 255 -17
rect 257 -19 260 -17
rect 253 -21 260 -19
rect 262 -15 268 -12
rect 284 -15 289 -8
rect 304 -8 311 -2
rect 388 0 394 2
rect 388 -2 390 0
rect 392 -2 394 0
rect 388 -4 394 -2
rect 409 0 416 2
rect 409 -2 411 0
rect 413 -2 416 0
rect 372 -7 377 -4
rect 304 -10 313 -8
rect 262 -21 270 -15
rect 272 -17 280 -15
rect 272 -19 275 -17
rect 277 -19 280 -17
rect 272 -21 280 -19
rect 282 -21 289 -15
rect 293 -12 300 -10
rect 293 -14 295 -12
rect 297 -14 300 -12
rect 293 -16 300 -14
rect 295 -19 300 -16
rect 302 -19 313 -10
rect 315 -19 320 -8
rect 322 -10 329 -8
rect 322 -12 325 -10
rect 327 -12 329 -10
rect 348 -9 357 -7
rect 348 -11 350 -9
rect 352 -11 357 -9
rect 348 -12 357 -11
rect 322 -14 329 -12
rect 322 -19 327 -14
rect 336 -15 341 -12
rect 334 -17 341 -15
rect 334 -19 336 -17
rect 338 -19 341 -17
rect 334 -21 341 -19
rect 343 -16 357 -12
rect 359 -12 367 -7
rect 359 -14 362 -12
rect 364 -14 367 -12
rect 359 -16 367 -14
rect 369 -10 377 -7
rect 369 -12 372 -10
rect 374 -12 377 -10
rect 369 -16 377 -12
rect 379 -16 384 -4
rect 386 -16 394 -4
rect 409 -8 416 -2
rect 493 0 499 2
rect 493 -2 495 0
rect 497 -2 499 0
rect 493 -4 499 -2
rect 514 -4 520 -2
rect 477 -7 482 -4
rect 409 -10 418 -8
rect 398 -12 405 -10
rect 398 -14 400 -12
rect 402 -14 405 -12
rect 398 -16 405 -14
rect 343 -21 348 -16
rect 400 -19 405 -16
rect 407 -19 418 -10
rect 420 -19 425 -8
rect 427 -10 434 -8
rect 427 -12 430 -10
rect 432 -12 434 -10
rect 453 -9 462 -7
rect 453 -11 455 -9
rect 457 -11 462 -9
rect 453 -12 462 -11
rect 427 -14 434 -12
rect 427 -19 432 -14
rect 441 -15 446 -12
rect 439 -17 446 -15
rect 439 -19 441 -17
rect 443 -19 446 -17
rect 439 -21 446 -19
rect 448 -16 462 -12
rect 464 -12 472 -7
rect 464 -14 467 -12
rect 469 -14 472 -12
rect 464 -16 472 -14
rect 474 -10 482 -7
rect 474 -12 477 -10
rect 479 -12 482 -10
rect 474 -16 482 -12
rect 484 -16 489 -4
rect 491 -16 499 -4
rect 514 -6 516 -4
rect 518 -6 520 -4
rect 514 -8 520 -6
rect 533 -4 539 -2
rect 554 0 561 2
rect 554 -2 556 0
rect 558 -2 561 0
rect 533 -6 535 -4
rect 537 -6 539 -4
rect 533 -8 539 -6
rect 514 -12 518 -8
rect 505 -15 510 -12
rect 448 -21 453 -16
rect 503 -17 510 -15
rect 503 -19 505 -17
rect 507 -19 510 -17
rect 503 -21 510 -19
rect 512 -15 518 -12
rect 534 -15 539 -8
rect 554 -8 561 -2
rect 638 0 644 2
rect 638 -2 640 0
rect 642 -2 644 0
rect 638 -4 644 -2
rect 659 0 666 2
rect 659 -2 661 0
rect 663 -2 666 0
rect 622 -7 627 -4
rect 554 -10 563 -8
rect 512 -21 520 -15
rect 522 -17 530 -15
rect 522 -19 525 -17
rect 527 -19 530 -17
rect 522 -21 530 -19
rect 532 -21 539 -15
rect 543 -12 550 -10
rect 543 -14 545 -12
rect 547 -14 550 -12
rect 543 -16 550 -14
rect 545 -19 550 -16
rect 552 -19 563 -10
rect 565 -19 570 -8
rect 572 -10 579 -8
rect 572 -12 575 -10
rect 577 -12 579 -10
rect 598 -9 607 -7
rect 598 -11 600 -9
rect 602 -11 607 -9
rect 598 -12 607 -11
rect 572 -14 579 -12
rect 572 -19 577 -14
rect 586 -15 591 -12
rect 584 -17 591 -15
rect 584 -19 586 -17
rect 588 -19 591 -17
rect 584 -21 591 -19
rect 593 -16 607 -12
rect 609 -12 617 -7
rect 609 -14 612 -12
rect 614 -14 617 -12
rect 609 -16 617 -14
rect 619 -10 627 -7
rect 619 -12 622 -10
rect 624 -12 627 -10
rect 619 -16 627 -12
rect 629 -16 634 -4
rect 636 -16 644 -4
rect 659 -8 666 -2
rect 743 0 749 2
rect 743 -2 745 0
rect 747 -2 749 0
rect 743 -4 749 -2
rect 727 -7 732 -4
rect 659 -10 668 -8
rect 648 -12 655 -10
rect 648 -14 650 -12
rect 652 -14 655 -12
rect 648 -16 655 -14
rect 593 -21 598 -16
rect 650 -19 655 -16
rect 657 -19 668 -10
rect 670 -19 675 -8
rect 677 -10 684 -8
rect 677 -12 680 -10
rect 682 -12 684 -10
rect 703 -9 712 -7
rect 703 -11 705 -9
rect 707 -11 712 -9
rect 703 -12 712 -11
rect 677 -14 684 -12
rect 677 -19 682 -14
rect 691 -15 696 -12
rect 689 -17 696 -15
rect 689 -19 691 -17
rect 693 -19 696 -17
rect 689 -21 696 -19
rect 698 -16 712 -12
rect 714 -12 722 -7
rect 714 -14 717 -12
rect 719 -14 722 -12
rect 714 -16 722 -14
rect 724 -10 732 -7
rect 724 -12 727 -10
rect 729 -12 732 -10
rect 724 -16 732 -12
rect 734 -16 739 -4
rect 741 -16 749 -4
rect 698 -21 703 -16
<< pdif >>
rect 40 103 46 110
rect 19 94 26 103
rect 19 92 21 94
rect 23 92 26 94
rect 19 90 26 92
rect 28 101 36 103
rect 28 99 31 101
rect 33 99 36 101
rect 28 94 36 99
rect 28 92 31 94
rect 33 92 36 94
rect 28 90 36 92
rect 38 96 46 103
rect 38 94 41 96
rect 43 94 46 96
rect 38 92 46 94
rect 48 108 55 110
rect 48 106 51 108
rect 53 106 55 108
rect 48 101 55 106
rect 80 103 86 110
rect 48 99 51 101
rect 53 99 55 101
rect 48 97 55 99
rect 48 92 53 97
rect 59 94 66 103
rect 59 92 61 94
rect 63 92 66 94
rect 38 90 44 92
rect 59 90 66 92
rect 68 101 76 103
rect 68 99 71 101
rect 73 99 76 101
rect 68 94 76 99
rect 68 92 71 94
rect 73 92 76 94
rect 68 90 76 92
rect 78 96 86 103
rect 78 94 81 96
rect 83 94 86 96
rect 78 92 86 94
rect 88 108 95 110
rect 88 106 91 108
rect 93 106 95 108
rect 88 101 95 106
rect 88 99 91 101
rect 93 99 95 101
rect 88 97 95 99
rect 88 92 93 97
rect 108 95 113 110
rect 106 93 113 95
rect 78 90 84 92
rect 106 91 108 93
rect 110 91 113 93
rect 106 89 113 91
rect 108 83 113 89
rect 115 101 123 110
rect 115 99 118 101
rect 120 99 123 101
rect 115 92 123 99
rect 125 108 133 110
rect 125 106 128 108
rect 130 106 133 108
rect 125 101 133 106
rect 125 99 128 101
rect 130 99 133 101
rect 125 92 133 99
rect 135 94 149 110
rect 135 92 144 94
rect 146 92 149 94
rect 115 83 120 92
rect 137 87 149 92
rect 137 85 144 87
rect 146 85 149 87
rect 137 83 149 85
rect 151 108 158 110
rect 151 106 154 108
rect 156 106 158 108
rect 151 104 158 106
rect 151 83 156 104
rect 192 103 198 110
rect 171 94 178 103
rect 171 92 173 94
rect 175 92 178 94
rect 171 90 178 92
rect 180 101 188 103
rect 180 99 183 101
rect 185 99 188 101
rect 180 94 188 99
rect 180 92 183 94
rect 185 92 188 94
rect 180 90 188 92
rect 190 96 198 103
rect 190 94 193 96
rect 195 94 198 96
rect 190 92 198 94
rect 200 108 207 110
rect 200 106 203 108
rect 205 106 207 108
rect 200 101 207 106
rect 245 103 251 110
rect 200 99 203 101
rect 205 99 207 101
rect 200 97 207 99
rect 200 92 205 97
rect 224 94 231 103
rect 224 92 226 94
rect 228 92 231 94
rect 190 90 196 92
rect 224 90 231 92
rect 233 101 241 103
rect 233 99 236 101
rect 238 99 241 101
rect 233 94 241 99
rect 233 92 236 94
rect 238 92 241 94
rect 233 90 241 92
rect 243 96 251 103
rect 243 94 246 96
rect 248 94 251 96
rect 243 92 251 94
rect 253 108 260 110
rect 253 106 256 108
rect 258 106 260 108
rect 253 101 260 106
rect 285 103 291 110
rect 253 99 256 101
rect 258 99 260 101
rect 253 97 260 99
rect 253 92 258 97
rect 264 94 271 103
rect 264 92 266 94
rect 268 92 271 94
rect 243 90 249 92
rect 264 90 271 92
rect 273 101 281 103
rect 273 99 276 101
rect 278 99 281 101
rect 273 94 281 99
rect 273 92 276 94
rect 278 92 281 94
rect 273 90 281 92
rect 283 96 291 103
rect 283 94 286 96
rect 288 94 291 96
rect 283 92 291 94
rect 293 108 300 110
rect 293 106 296 108
rect 298 106 300 108
rect 293 101 300 106
rect 293 99 296 101
rect 298 99 300 101
rect 293 97 300 99
rect 293 92 298 97
rect 313 95 318 110
rect 311 93 318 95
rect 283 90 289 92
rect 311 91 313 93
rect 315 91 318 93
rect 311 89 318 91
rect 313 83 318 89
rect 320 101 328 110
rect 320 99 323 101
rect 325 99 328 101
rect 320 92 328 99
rect 330 108 338 110
rect 330 106 333 108
rect 335 106 338 108
rect 330 101 338 106
rect 330 99 333 101
rect 335 99 338 101
rect 330 92 338 99
rect 340 94 354 110
rect 340 92 349 94
rect 351 92 354 94
rect 320 83 325 92
rect 342 87 354 92
rect 342 85 349 87
rect 351 85 354 87
rect 342 83 354 85
rect 356 108 363 110
rect 356 106 359 108
rect 361 106 363 108
rect 356 104 363 106
rect 356 83 361 104
rect 397 103 403 110
rect 376 94 383 103
rect 376 92 378 94
rect 380 92 383 94
rect 376 90 383 92
rect 385 101 393 103
rect 385 99 388 101
rect 390 99 393 101
rect 385 94 393 99
rect 385 92 388 94
rect 390 92 393 94
rect 385 90 393 92
rect 395 96 403 103
rect 395 94 398 96
rect 400 94 403 96
rect 395 92 403 94
rect 405 108 412 110
rect 405 106 408 108
rect 410 106 412 108
rect 405 101 412 106
rect 405 99 408 101
rect 410 99 412 101
rect 405 97 412 99
rect 405 92 410 97
rect 395 90 401 92
rect 30 62 36 64
rect 21 57 26 62
rect 19 55 26 57
rect 19 53 21 55
rect 23 53 26 55
rect 19 48 26 53
rect 19 46 21 48
rect 23 46 26 48
rect 19 44 26 46
rect 28 60 36 62
rect 28 58 31 60
rect 33 58 36 60
rect 28 51 36 58
rect 38 62 46 64
rect 38 60 41 62
rect 43 60 46 62
rect 38 55 46 60
rect 38 53 41 55
rect 43 53 46 55
rect 38 51 46 53
rect 48 62 55 64
rect 48 60 51 62
rect 53 60 55 62
rect 48 51 55 60
rect 59 62 66 64
rect 59 60 61 62
rect 63 60 66 62
rect 59 51 66 60
rect 68 62 76 64
rect 68 60 71 62
rect 73 60 76 62
rect 68 55 76 60
rect 68 53 71 55
rect 73 53 76 55
rect 68 51 76 53
rect 78 62 84 64
rect 110 62 116 64
rect 78 60 86 62
rect 78 58 81 60
rect 83 58 86 60
rect 78 51 86 58
rect 28 44 34 51
rect 80 44 86 51
rect 88 57 93 62
rect 101 57 106 62
rect 88 55 95 57
rect 88 53 91 55
rect 93 53 95 55
rect 88 48 95 53
rect 88 46 91 48
rect 93 46 95 48
rect 88 44 95 46
rect 99 55 106 57
rect 99 53 101 55
rect 103 53 106 55
rect 99 48 106 53
rect 99 46 101 48
rect 103 46 106 48
rect 99 44 106 46
rect 108 60 116 62
rect 108 58 111 60
rect 113 58 116 60
rect 108 51 116 58
rect 118 62 126 64
rect 118 60 121 62
rect 123 60 126 62
rect 118 55 126 60
rect 118 53 121 55
rect 123 53 126 55
rect 118 51 126 53
rect 128 62 135 64
rect 128 60 131 62
rect 133 60 135 62
rect 128 51 135 60
rect 108 44 114 51
rect 150 50 155 71
rect 148 48 155 50
rect 148 46 150 48
rect 152 46 155 48
rect 148 44 155 46
rect 157 69 169 71
rect 157 67 160 69
rect 162 67 169 69
rect 157 62 169 67
rect 186 62 191 71
rect 157 60 160 62
rect 162 60 171 62
rect 157 44 171 60
rect 173 55 181 62
rect 173 53 176 55
rect 178 53 181 55
rect 173 48 181 53
rect 173 46 176 48
rect 178 46 181 48
rect 173 44 181 46
rect 183 55 191 62
rect 183 53 186 55
rect 188 53 191 55
rect 183 44 191 53
rect 193 65 198 71
rect 193 63 200 65
rect 193 61 196 63
rect 198 61 200 63
rect 235 62 241 64
rect 193 59 200 61
rect 193 44 198 59
rect 226 57 231 62
rect 224 55 231 57
rect 224 53 226 55
rect 228 53 231 55
rect 224 48 231 53
rect 224 46 226 48
rect 228 46 231 48
rect 224 44 231 46
rect 233 60 241 62
rect 233 58 236 60
rect 238 58 241 60
rect 233 51 241 58
rect 243 62 251 64
rect 243 60 246 62
rect 248 60 251 62
rect 243 55 251 60
rect 243 53 246 55
rect 248 53 251 55
rect 243 51 251 53
rect 253 62 260 64
rect 253 60 256 62
rect 258 60 260 62
rect 253 51 260 60
rect 264 62 271 64
rect 264 60 266 62
rect 268 60 271 62
rect 264 51 271 60
rect 273 62 281 64
rect 273 60 276 62
rect 278 60 281 62
rect 273 55 281 60
rect 273 53 276 55
rect 278 53 281 55
rect 273 51 281 53
rect 283 62 289 64
rect 315 62 321 64
rect 283 60 291 62
rect 283 58 286 60
rect 288 58 291 60
rect 283 51 291 58
rect 233 44 239 51
rect 285 44 291 51
rect 293 57 298 62
rect 306 57 311 62
rect 293 55 300 57
rect 293 53 296 55
rect 298 53 300 55
rect 293 48 300 53
rect 293 46 296 48
rect 298 46 300 48
rect 293 44 300 46
rect 304 55 311 57
rect 304 53 306 55
rect 308 53 311 55
rect 304 48 311 53
rect 304 46 306 48
rect 308 46 311 48
rect 304 44 311 46
rect 313 60 321 62
rect 313 58 316 60
rect 318 58 321 60
rect 313 51 321 58
rect 323 62 331 64
rect 323 60 326 62
rect 328 60 331 62
rect 323 55 331 60
rect 323 53 326 55
rect 328 53 331 55
rect 323 51 331 53
rect 333 62 340 64
rect 333 60 336 62
rect 338 60 340 62
rect 333 51 340 60
rect 313 44 319 51
rect 355 50 360 71
rect 353 48 360 50
rect 353 46 355 48
rect 357 46 360 48
rect 353 44 360 46
rect 362 69 374 71
rect 362 67 365 69
rect 367 67 374 69
rect 362 62 374 67
rect 391 62 396 71
rect 362 60 365 62
rect 367 60 376 62
rect 362 44 376 60
rect 378 55 386 62
rect 378 53 381 55
rect 383 53 386 55
rect 378 48 386 53
rect 378 46 381 48
rect 383 46 386 48
rect 378 44 386 46
rect 388 55 396 62
rect 388 53 391 55
rect 393 53 396 55
rect 388 44 396 53
rect 398 65 403 71
rect 398 63 405 65
rect 398 61 401 63
rect 403 61 405 63
rect 398 59 405 61
rect 398 44 403 59
rect -245 -38 -240 -33
rect -247 -40 -240 -38
rect -247 -42 -245 -40
rect -243 -42 -240 -40
rect -247 -47 -240 -42
rect -247 -49 -245 -47
rect -243 -49 -240 -47
rect -247 -51 -240 -49
rect -238 -40 -230 -33
rect -207 -36 -200 -34
rect -207 -38 -205 -36
rect -203 -38 -200 -36
rect -238 -51 -227 -40
rect -236 -57 -227 -51
rect -236 -59 -234 -57
rect -232 -59 -227 -57
rect -236 -61 -227 -59
rect -225 -61 -220 -40
rect -218 -48 -213 -40
rect -207 -43 -200 -38
rect -207 -45 -205 -43
rect -203 -45 -200 -43
rect -207 -47 -200 -45
rect -218 -50 -211 -48
rect -218 -52 -215 -50
rect -213 -52 -211 -50
rect -205 -52 -200 -47
rect -198 -41 -192 -34
rect -158 -36 -151 -34
rect -158 -38 -156 -36
rect -154 -38 -151 -36
rect -158 -40 -151 -38
rect -198 -48 -190 -41
rect -198 -50 -195 -48
rect -193 -50 -190 -48
rect -198 -52 -190 -50
rect -218 -54 -211 -52
rect -218 -61 -213 -54
rect -196 -54 -190 -52
rect -188 -43 -180 -41
rect -188 -45 -185 -43
rect -183 -45 -180 -43
rect -188 -50 -180 -45
rect -188 -52 -185 -50
rect -183 -52 -180 -50
rect -188 -54 -180 -52
rect -178 -50 -171 -41
rect -178 -52 -175 -50
rect -173 -52 -171 -50
rect -178 -54 -171 -52
rect -156 -61 -151 -40
rect -149 -50 -135 -34
rect -149 -52 -146 -50
rect -144 -52 -135 -50
rect -133 -36 -125 -34
rect -133 -38 -130 -36
rect -128 -38 -125 -36
rect -133 -43 -125 -38
rect -133 -45 -130 -43
rect -128 -45 -125 -43
rect -133 -52 -125 -45
rect -123 -43 -115 -34
rect -123 -45 -120 -43
rect -118 -45 -115 -43
rect -123 -52 -115 -45
rect -149 -57 -137 -52
rect -149 -59 -146 -57
rect -144 -59 -137 -57
rect -149 -61 -137 -59
rect -120 -61 -115 -52
rect -113 -49 -108 -34
rect -102 -36 -95 -34
rect -102 -38 -100 -36
rect -98 -38 -95 -36
rect -102 -43 -95 -38
rect -102 -45 -100 -43
rect -98 -45 -95 -43
rect -102 -47 -95 -45
rect -113 -51 -106 -49
rect -113 -53 -110 -51
rect -108 -53 -106 -51
rect -100 -52 -95 -47
rect -93 -41 -87 -34
rect -53 -36 -46 -34
rect -53 -38 -51 -36
rect -49 -38 -46 -36
rect -53 -40 -46 -38
rect -93 -48 -85 -41
rect -93 -50 -90 -48
rect -88 -50 -85 -48
rect -93 -52 -85 -50
rect -113 -55 -106 -53
rect -113 -61 -108 -55
rect -91 -54 -85 -52
rect -83 -43 -75 -41
rect -83 -45 -80 -43
rect -78 -45 -75 -43
rect -83 -50 -75 -45
rect -83 -52 -80 -50
rect -78 -52 -75 -50
rect -83 -54 -75 -52
rect -73 -50 -66 -41
rect -73 -52 -70 -50
rect -68 -52 -66 -50
rect -73 -54 -66 -52
rect -51 -61 -46 -40
rect -44 -50 -30 -34
rect -44 -52 -41 -50
rect -39 -52 -30 -50
rect -28 -36 -20 -34
rect -28 -38 -25 -36
rect -23 -38 -20 -36
rect -28 -43 -20 -38
rect -28 -45 -25 -43
rect -23 -45 -20 -43
rect -28 -52 -20 -45
rect -18 -43 -10 -34
rect -18 -45 -15 -43
rect -13 -45 -10 -43
rect -18 -52 -10 -45
rect -44 -57 -32 -52
rect -44 -59 -41 -57
rect -39 -59 -32 -57
rect -44 -61 -32 -59
rect -15 -61 -10 -52
rect -8 -49 -3 -34
rect 5 -38 10 -33
rect 3 -40 10 -38
rect 3 -42 5 -40
rect 7 -42 10 -40
rect 3 -47 10 -42
rect 3 -49 5 -47
rect 7 -49 10 -47
rect -8 -51 -1 -49
rect 3 -51 10 -49
rect 12 -40 20 -33
rect 43 -36 50 -34
rect 43 -38 45 -36
rect 47 -38 50 -36
rect 12 -51 23 -40
rect -8 -53 -5 -51
rect -3 -53 -1 -51
rect -8 -55 -1 -53
rect -8 -61 -3 -55
rect 14 -57 23 -51
rect 14 -59 16 -57
rect 18 -59 23 -57
rect 14 -61 23 -59
rect 25 -61 30 -40
rect 32 -48 37 -40
rect 43 -43 50 -38
rect 43 -45 45 -43
rect 47 -45 50 -43
rect 43 -47 50 -45
rect 32 -50 39 -48
rect 32 -52 35 -50
rect 37 -52 39 -50
rect 45 -52 50 -47
rect 52 -41 58 -34
rect 92 -36 99 -34
rect 92 -38 94 -36
rect 96 -38 99 -36
rect 92 -40 99 -38
rect 52 -48 60 -41
rect 52 -50 55 -48
rect 57 -50 60 -48
rect 52 -52 60 -50
rect 32 -54 39 -52
rect 32 -61 37 -54
rect 54 -54 60 -52
rect 62 -43 70 -41
rect 62 -45 65 -43
rect 67 -45 70 -43
rect 62 -50 70 -45
rect 62 -52 65 -50
rect 67 -52 70 -50
rect 62 -54 70 -52
rect 72 -50 79 -41
rect 72 -52 75 -50
rect 77 -52 79 -50
rect 72 -54 79 -52
rect 94 -61 99 -40
rect 101 -50 115 -34
rect 101 -52 104 -50
rect 106 -52 115 -50
rect 117 -36 125 -34
rect 117 -38 120 -36
rect 122 -38 125 -36
rect 117 -43 125 -38
rect 117 -45 120 -43
rect 122 -45 125 -43
rect 117 -52 125 -45
rect 127 -43 135 -34
rect 127 -45 130 -43
rect 132 -45 135 -43
rect 127 -52 135 -45
rect 101 -57 113 -52
rect 101 -59 104 -57
rect 106 -59 113 -57
rect 101 -61 113 -59
rect 130 -61 135 -52
rect 137 -49 142 -34
rect 148 -36 155 -34
rect 148 -38 150 -36
rect 152 -38 155 -36
rect 148 -43 155 -38
rect 148 -45 150 -43
rect 152 -45 155 -43
rect 148 -47 155 -45
rect 137 -51 144 -49
rect 137 -53 140 -51
rect 142 -53 144 -51
rect 150 -52 155 -47
rect 157 -41 163 -34
rect 197 -36 204 -34
rect 197 -38 199 -36
rect 201 -38 204 -36
rect 197 -40 204 -38
rect 157 -48 165 -41
rect 157 -50 160 -48
rect 162 -50 165 -48
rect 157 -52 165 -50
rect 137 -55 144 -53
rect 137 -61 142 -55
rect 159 -54 165 -52
rect 167 -43 175 -41
rect 167 -45 170 -43
rect 172 -45 175 -43
rect 167 -50 175 -45
rect 167 -52 170 -50
rect 172 -52 175 -50
rect 167 -54 175 -52
rect 177 -50 184 -41
rect 177 -52 180 -50
rect 182 -52 184 -50
rect 177 -54 184 -52
rect 199 -61 204 -40
rect 206 -50 220 -34
rect 206 -52 209 -50
rect 211 -52 220 -50
rect 222 -36 230 -34
rect 222 -38 225 -36
rect 227 -38 230 -36
rect 222 -43 230 -38
rect 222 -45 225 -43
rect 227 -45 230 -43
rect 222 -52 230 -45
rect 232 -43 240 -34
rect 232 -45 235 -43
rect 237 -45 240 -43
rect 232 -52 240 -45
rect 206 -57 218 -52
rect 206 -59 209 -57
rect 211 -59 218 -57
rect 206 -61 218 -59
rect 235 -61 240 -52
rect 242 -49 247 -34
rect 255 -38 260 -33
rect 253 -40 260 -38
rect 253 -42 255 -40
rect 257 -42 260 -40
rect 253 -47 260 -42
rect 253 -49 255 -47
rect 257 -49 260 -47
rect 242 -51 249 -49
rect 253 -51 260 -49
rect 262 -40 270 -33
rect 293 -36 300 -34
rect 293 -38 295 -36
rect 297 -38 300 -36
rect 262 -51 273 -40
rect 242 -53 245 -51
rect 247 -53 249 -51
rect 242 -55 249 -53
rect 242 -61 247 -55
rect 264 -57 273 -51
rect 264 -59 266 -57
rect 268 -59 273 -57
rect 264 -61 273 -59
rect 275 -61 280 -40
rect 282 -48 287 -40
rect 293 -43 300 -38
rect 293 -45 295 -43
rect 297 -45 300 -43
rect 293 -47 300 -45
rect 282 -50 289 -48
rect 282 -52 285 -50
rect 287 -52 289 -50
rect 295 -52 300 -47
rect 302 -41 308 -34
rect 342 -36 349 -34
rect 342 -38 344 -36
rect 346 -38 349 -36
rect 342 -40 349 -38
rect 302 -48 310 -41
rect 302 -50 305 -48
rect 307 -50 310 -48
rect 302 -52 310 -50
rect 282 -54 289 -52
rect 282 -61 287 -54
rect 304 -54 310 -52
rect 312 -43 320 -41
rect 312 -45 315 -43
rect 317 -45 320 -43
rect 312 -50 320 -45
rect 312 -52 315 -50
rect 317 -52 320 -50
rect 312 -54 320 -52
rect 322 -50 329 -41
rect 322 -52 325 -50
rect 327 -52 329 -50
rect 322 -54 329 -52
rect 344 -61 349 -40
rect 351 -50 365 -34
rect 351 -52 354 -50
rect 356 -52 365 -50
rect 367 -36 375 -34
rect 367 -38 370 -36
rect 372 -38 375 -36
rect 367 -43 375 -38
rect 367 -45 370 -43
rect 372 -45 375 -43
rect 367 -52 375 -45
rect 377 -43 385 -34
rect 377 -45 380 -43
rect 382 -45 385 -43
rect 377 -52 385 -45
rect 351 -57 363 -52
rect 351 -59 354 -57
rect 356 -59 363 -57
rect 351 -61 363 -59
rect 380 -61 385 -52
rect 387 -49 392 -34
rect 398 -36 405 -34
rect 398 -38 400 -36
rect 402 -38 405 -36
rect 398 -43 405 -38
rect 398 -45 400 -43
rect 402 -45 405 -43
rect 398 -47 405 -45
rect 387 -51 394 -49
rect 387 -53 390 -51
rect 392 -53 394 -51
rect 400 -52 405 -47
rect 407 -41 413 -34
rect 447 -36 454 -34
rect 447 -38 449 -36
rect 451 -38 454 -36
rect 447 -40 454 -38
rect 407 -48 415 -41
rect 407 -50 410 -48
rect 412 -50 415 -48
rect 407 -52 415 -50
rect 387 -55 394 -53
rect 387 -61 392 -55
rect 409 -54 415 -52
rect 417 -43 425 -41
rect 417 -45 420 -43
rect 422 -45 425 -43
rect 417 -50 425 -45
rect 417 -52 420 -50
rect 422 -52 425 -50
rect 417 -54 425 -52
rect 427 -50 434 -41
rect 427 -52 430 -50
rect 432 -52 434 -50
rect 427 -54 434 -52
rect 449 -61 454 -40
rect 456 -50 470 -34
rect 456 -52 459 -50
rect 461 -52 470 -50
rect 472 -36 480 -34
rect 472 -38 475 -36
rect 477 -38 480 -36
rect 472 -43 480 -38
rect 472 -45 475 -43
rect 477 -45 480 -43
rect 472 -52 480 -45
rect 482 -43 490 -34
rect 482 -45 485 -43
rect 487 -45 490 -43
rect 482 -52 490 -45
rect 456 -57 468 -52
rect 456 -59 459 -57
rect 461 -59 468 -57
rect 456 -61 468 -59
rect 485 -61 490 -52
rect 492 -49 497 -34
rect 505 -38 510 -33
rect 503 -40 510 -38
rect 503 -42 505 -40
rect 507 -42 510 -40
rect 503 -47 510 -42
rect 503 -49 505 -47
rect 507 -49 510 -47
rect 492 -51 499 -49
rect 503 -51 510 -49
rect 512 -40 520 -33
rect 543 -36 550 -34
rect 543 -38 545 -36
rect 547 -38 550 -36
rect 512 -51 523 -40
rect 492 -53 495 -51
rect 497 -53 499 -51
rect 492 -55 499 -53
rect 492 -61 497 -55
rect 514 -57 523 -51
rect 514 -59 516 -57
rect 518 -59 523 -57
rect 514 -61 523 -59
rect 525 -61 530 -40
rect 532 -48 537 -40
rect 543 -43 550 -38
rect 543 -45 545 -43
rect 547 -45 550 -43
rect 543 -47 550 -45
rect 532 -50 539 -48
rect 532 -52 535 -50
rect 537 -52 539 -50
rect 545 -52 550 -47
rect 552 -41 558 -34
rect 592 -36 599 -34
rect 592 -38 594 -36
rect 596 -38 599 -36
rect 592 -40 599 -38
rect 552 -48 560 -41
rect 552 -50 555 -48
rect 557 -50 560 -48
rect 552 -52 560 -50
rect 532 -54 539 -52
rect 532 -61 537 -54
rect 554 -54 560 -52
rect 562 -43 570 -41
rect 562 -45 565 -43
rect 567 -45 570 -43
rect 562 -50 570 -45
rect 562 -52 565 -50
rect 567 -52 570 -50
rect 562 -54 570 -52
rect 572 -50 579 -41
rect 572 -52 575 -50
rect 577 -52 579 -50
rect 572 -54 579 -52
rect 594 -61 599 -40
rect 601 -50 615 -34
rect 601 -52 604 -50
rect 606 -52 615 -50
rect 617 -36 625 -34
rect 617 -38 620 -36
rect 622 -38 625 -36
rect 617 -43 625 -38
rect 617 -45 620 -43
rect 622 -45 625 -43
rect 617 -52 625 -45
rect 627 -43 635 -34
rect 627 -45 630 -43
rect 632 -45 635 -43
rect 627 -52 635 -45
rect 601 -57 613 -52
rect 601 -59 604 -57
rect 606 -59 613 -57
rect 601 -61 613 -59
rect 630 -61 635 -52
rect 637 -49 642 -34
rect 648 -36 655 -34
rect 648 -38 650 -36
rect 652 -38 655 -36
rect 648 -43 655 -38
rect 648 -45 650 -43
rect 652 -45 655 -43
rect 648 -47 655 -45
rect 637 -51 644 -49
rect 637 -53 640 -51
rect 642 -53 644 -51
rect 650 -52 655 -47
rect 657 -41 663 -34
rect 697 -36 704 -34
rect 697 -38 699 -36
rect 701 -38 704 -36
rect 697 -40 704 -38
rect 657 -48 665 -41
rect 657 -50 660 -48
rect 662 -50 665 -48
rect 657 -52 665 -50
rect 637 -55 644 -53
rect 637 -61 642 -55
rect 659 -54 665 -52
rect 667 -43 675 -41
rect 667 -45 670 -43
rect 672 -45 675 -43
rect 667 -50 675 -45
rect 667 -52 670 -50
rect 672 -52 675 -50
rect 667 -54 675 -52
rect 677 -50 684 -41
rect 677 -52 680 -50
rect 682 -52 684 -50
rect 677 -54 684 -52
rect 699 -61 704 -40
rect 706 -50 720 -34
rect 706 -52 709 -50
rect 711 -52 720 -50
rect 722 -36 730 -34
rect 722 -38 725 -36
rect 727 -38 730 -36
rect 722 -43 730 -38
rect 722 -45 725 -43
rect 727 -45 730 -43
rect 722 -52 730 -45
rect 732 -43 740 -34
rect 732 -45 735 -43
rect 737 -45 740 -43
rect 732 -52 740 -45
rect 706 -57 718 -52
rect 706 -59 709 -57
rect 711 -59 718 -57
rect 706 -61 718 -59
rect 735 -61 740 -52
rect 742 -49 747 -34
rect 742 -51 749 -49
rect 742 -53 745 -51
rect 747 -53 749 -51
rect 742 -55 749 -53
rect 742 -61 747 -55
<< alu1 >>
rect 9 144 412 149
rect 9 142 40 144
rect 42 142 50 144
rect 52 142 80 144
rect 82 142 90 144
rect 92 142 108 144
rect 110 142 161 144
rect 163 142 192 144
rect 194 142 202 144
rect 204 142 245 144
rect 247 142 255 144
rect 257 142 285 144
rect 287 142 295 144
rect 297 142 313 144
rect 315 142 366 144
rect 368 142 397 144
rect 399 142 407 144
rect 409 142 412 144
rect 9 141 412 142
rect 26 119 31 128
rect 43 132 55 136
rect 43 130 51 132
rect 53 130 55 132
rect 51 127 55 130
rect 26 118 40 119
rect 26 116 34 118
rect 36 116 37 118
rect 39 116 40 118
rect 26 115 40 116
rect 19 110 32 111
rect 19 108 24 110
rect 26 108 32 110
rect 19 107 32 108
rect 19 102 23 107
rect 51 125 52 127
rect 54 125 55 127
rect 51 110 55 125
rect 66 119 71 128
rect 83 132 95 136
rect 83 130 91 132
rect 93 130 95 132
rect 66 118 80 119
rect 66 116 74 118
rect 76 116 77 118
rect 79 116 80 118
rect 66 115 80 116
rect 19 100 20 102
rect 22 100 23 102
rect 19 98 23 100
rect 50 108 55 110
rect 50 106 51 108
rect 53 106 55 108
rect 50 101 55 106
rect 50 99 51 101
rect 53 99 55 101
rect 50 97 55 99
rect 59 110 72 111
rect 59 108 64 110
rect 66 108 72 110
rect 59 107 72 108
rect 59 103 63 107
rect 91 110 95 130
rect 59 101 60 103
rect 62 101 63 103
rect 59 98 63 101
rect 90 108 95 110
rect 90 106 91 108
rect 93 106 95 108
rect 90 104 95 106
rect 90 102 91 104
rect 93 102 95 104
rect 90 101 95 102
rect 90 99 91 101
rect 93 99 95 101
rect 90 97 95 99
rect 106 134 130 135
rect 106 132 126 134
rect 128 132 130 134
rect 106 131 130 132
rect 106 103 110 131
rect 145 127 158 128
rect 145 125 153 127
rect 155 125 158 127
rect 145 123 158 125
rect 145 121 146 123
rect 148 122 158 123
rect 148 121 150 122
rect 106 101 122 103
rect 106 99 118 101
rect 120 99 122 101
rect 106 98 122 99
rect 145 114 150 121
rect 178 127 183 128
rect 178 125 180 127
rect 182 125 183 127
rect 178 119 183 125
rect 195 132 207 136
rect 195 130 203 132
rect 205 130 207 132
rect 178 118 192 119
rect 178 116 186 118
rect 188 116 192 118
rect 178 115 192 116
rect 161 111 166 112
rect 161 110 167 111
rect 171 110 184 111
rect 161 108 162 110
rect 164 108 176 110
rect 178 108 184 110
rect 161 107 184 108
rect 161 105 175 107
rect 161 96 166 105
rect 171 104 175 105
rect 203 115 207 130
rect 231 119 236 128
rect 248 132 260 136
rect 248 130 256 132
rect 258 130 260 132
rect 256 127 260 130
rect 231 118 245 119
rect 231 116 239 118
rect 241 116 242 118
rect 244 116 245 118
rect 231 115 245 116
rect 203 113 204 115
rect 206 113 207 115
rect 203 110 207 113
rect 171 102 172 104
rect 174 102 175 104
rect 171 98 175 102
rect 202 108 207 110
rect 202 106 203 108
rect 205 106 207 108
rect 202 101 207 106
rect 154 90 166 96
rect 202 99 203 101
rect 205 99 207 101
rect 202 97 207 99
rect 224 110 237 111
rect 224 108 229 110
rect 231 108 237 110
rect 224 107 237 108
rect 224 102 228 107
rect 256 125 257 127
rect 259 125 260 127
rect 256 110 260 125
rect 271 119 276 128
rect 288 132 300 136
rect 288 130 296 132
rect 298 130 300 132
rect 271 118 285 119
rect 271 116 279 118
rect 281 116 282 118
rect 284 116 285 118
rect 271 115 285 116
rect 224 100 225 102
rect 227 100 228 102
rect 224 98 228 100
rect 255 108 260 110
rect 255 106 256 108
rect 258 106 260 108
rect 255 101 260 106
rect 255 99 256 101
rect 258 99 260 101
rect 255 97 260 99
rect 264 110 277 111
rect 264 108 269 110
rect 271 108 277 110
rect 264 107 277 108
rect 264 103 268 107
rect 296 110 300 130
rect 264 101 265 103
rect 267 101 268 103
rect 264 98 268 101
rect 295 108 300 110
rect 295 106 296 108
rect 298 106 300 108
rect 295 104 300 106
rect 295 102 296 104
rect 298 102 300 104
rect 295 101 300 102
rect 295 99 296 101
rect 298 99 300 101
rect 295 97 300 99
rect 311 134 335 135
rect 311 132 331 134
rect 333 132 335 134
rect 311 131 335 132
rect 311 103 315 131
rect 350 127 363 128
rect 350 125 358 127
rect 360 125 363 127
rect 350 123 363 125
rect 350 121 351 123
rect 353 122 363 123
rect 353 121 355 122
rect 311 101 327 103
rect 311 99 323 101
rect 325 99 327 101
rect 311 98 327 99
rect 350 114 355 121
rect 383 127 388 128
rect 383 125 385 127
rect 387 125 388 127
rect 383 119 388 125
rect 400 132 412 136
rect 400 130 408 132
rect 410 130 412 132
rect 383 118 397 119
rect 383 116 391 118
rect 393 116 397 118
rect 383 115 397 116
rect 366 111 371 112
rect 366 110 372 111
rect 376 110 389 111
rect 366 108 367 110
rect 369 108 381 110
rect 383 108 389 110
rect 366 107 389 108
rect 366 105 380 107
rect 366 96 371 105
rect 376 104 380 105
rect 408 115 412 130
rect 408 113 409 115
rect 411 113 412 115
rect 408 110 412 113
rect 376 102 377 104
rect 379 102 380 104
rect 376 98 380 102
rect 407 108 412 110
rect 407 106 408 108
rect 410 106 412 108
rect 407 101 412 106
rect 359 90 371 96
rect 407 99 408 101
rect 410 99 412 101
rect 407 97 412 99
rect 18 84 412 85
rect 18 82 50 84
rect 52 82 90 84
rect 92 82 128 84
rect 130 82 202 84
rect 204 82 255 84
rect 257 82 295 84
rect 297 82 333 84
rect 335 82 407 84
rect 409 82 412 84
rect 18 72 412 82
rect 18 70 22 72
rect 24 70 90 72
rect 92 70 102 72
rect 104 70 176 72
rect 178 70 227 72
rect 229 70 295 72
rect 297 70 307 72
rect 309 70 381 72
rect 383 70 412 72
rect 18 69 412 70
rect 19 55 24 57
rect 19 53 21 55
rect 23 53 24 55
rect 19 48 24 53
rect 19 46 21 48
rect 23 46 24 48
rect 19 44 24 46
rect 51 55 55 56
rect 51 53 52 55
rect 54 53 55 55
rect 19 24 23 44
rect 51 47 55 53
rect 42 46 55 47
rect 42 44 48 46
rect 50 44 55 46
rect 42 43 55 44
rect 59 47 63 56
rect 90 55 95 57
rect 59 46 72 47
rect 59 44 60 46
rect 62 44 64 46
rect 66 44 72 46
rect 59 43 72 44
rect 34 38 48 39
rect 34 36 35 38
rect 37 36 38 38
rect 40 36 48 38
rect 34 35 48 36
rect 19 22 21 24
rect 23 22 31 24
rect 19 18 31 22
rect 43 26 48 35
rect 66 38 80 39
rect 66 36 74 38
rect 76 36 77 38
rect 79 36 80 38
rect 66 35 80 36
rect 90 53 91 55
rect 93 53 95 55
rect 90 48 95 53
rect 90 46 91 48
rect 93 46 95 48
rect 90 44 95 46
rect 66 26 71 35
rect 91 29 95 44
rect 91 27 92 29
rect 94 27 95 29
rect 91 24 95 27
rect 83 22 91 24
rect 93 22 95 24
rect 83 18 95 22
rect 99 55 104 57
rect 99 53 101 55
rect 103 53 104 55
rect 140 62 152 64
rect 140 60 148 62
rect 150 60 152 62
rect 140 58 152 60
rect 99 48 104 53
rect 99 46 101 48
rect 103 46 104 48
rect 99 44 104 46
rect 99 24 103 44
rect 131 49 135 56
rect 140 49 145 58
rect 131 47 145 49
rect 122 46 145 47
rect 122 44 128 46
rect 130 44 142 46
rect 144 44 145 46
rect 122 43 135 44
rect 139 43 145 44
rect 140 42 145 43
rect 114 38 128 39
rect 114 36 118 38
rect 120 36 128 38
rect 114 35 128 36
rect 99 22 101 24
rect 103 22 111 24
rect 99 18 111 22
rect 123 29 128 35
rect 123 27 124 29
rect 126 27 128 29
rect 123 26 128 27
rect 156 33 161 40
rect 184 55 200 56
rect 184 53 186 55
rect 188 53 200 55
rect 184 51 200 53
rect 156 32 158 33
rect 148 31 158 32
rect 160 31 161 33
rect 148 29 161 31
rect 148 27 151 29
rect 153 27 161 29
rect 148 26 161 27
rect 196 23 200 51
rect 176 22 200 23
rect 176 20 178 22
rect 180 20 200 22
rect 176 19 200 20
rect 224 55 229 57
rect 224 53 226 55
rect 228 53 229 55
rect 224 48 229 53
rect 224 46 226 48
rect 228 46 229 48
rect 224 44 229 46
rect 256 55 260 56
rect 256 53 257 55
rect 259 53 260 55
rect 224 24 228 44
rect 256 47 260 53
rect 247 46 260 47
rect 247 44 253 46
rect 255 44 260 46
rect 247 43 260 44
rect 264 47 268 56
rect 295 55 300 57
rect 264 46 277 47
rect 264 44 265 46
rect 267 44 269 46
rect 271 44 277 46
rect 264 43 277 44
rect 239 38 253 39
rect 239 36 240 38
rect 242 36 243 38
rect 245 36 253 38
rect 239 35 253 36
rect 224 22 226 24
rect 228 22 236 24
rect 224 18 236 22
rect 248 26 253 35
rect 271 38 285 39
rect 271 36 279 38
rect 281 36 282 38
rect 284 36 285 38
rect 271 35 285 36
rect 295 53 296 55
rect 298 53 300 55
rect 295 48 300 53
rect 295 46 296 48
rect 298 46 300 48
rect 295 44 300 46
rect 271 26 276 35
rect 296 29 300 44
rect 296 27 297 29
rect 299 27 300 29
rect 296 24 300 27
rect 288 22 296 24
rect 298 22 300 24
rect 288 18 300 22
rect 304 55 309 57
rect 304 53 306 55
rect 308 53 309 55
rect 345 62 357 64
rect 345 60 353 62
rect 355 60 357 62
rect 345 58 357 60
rect 304 48 309 53
rect 304 46 306 48
rect 308 46 309 48
rect 304 44 309 46
rect 304 24 308 44
rect 336 49 340 56
rect 345 49 350 58
rect 336 47 350 49
rect 327 46 350 47
rect 327 44 333 46
rect 335 44 347 46
rect 349 44 350 46
rect 327 43 340 44
rect 344 43 350 44
rect 345 42 350 43
rect 319 38 333 39
rect 319 36 323 38
rect 325 36 333 38
rect 319 35 333 36
rect 304 22 306 24
rect 308 22 316 24
rect 304 18 316 22
rect 328 29 333 35
rect 328 27 329 29
rect 331 27 333 29
rect 328 26 333 27
rect 361 33 366 40
rect 389 55 405 56
rect 389 53 391 55
rect 393 53 405 55
rect 389 51 405 53
rect 361 32 363 33
rect 353 31 363 32
rect 365 31 366 33
rect 353 29 366 31
rect 353 27 356 29
rect 358 27 366 29
rect 353 26 366 27
rect 401 23 405 51
rect 381 22 405 23
rect 381 20 383 22
rect 385 20 405 22
rect 381 19 405 20
rect 9 12 409 13
rect 9 10 22 12
rect 24 10 32 12
rect 34 10 80 12
rect 82 10 90 12
rect 92 10 102 12
rect 104 10 112 12
rect 114 10 143 12
rect 145 10 196 12
rect 198 10 227 12
rect 229 10 237 12
rect 239 10 285 12
rect 287 10 295 12
rect 297 10 307 12
rect 309 10 317 12
rect 319 10 348 12
rect 350 10 401 12
rect 403 10 409 12
rect 9 5 409 10
rect -251 0 753 5
rect -251 -2 -244 0
rect -242 -2 -204 0
rect -202 -2 -194 0
rect -192 -2 -163 0
rect -161 -2 -110 0
rect -108 -2 -99 0
rect -97 -2 -89 0
rect -87 -2 -58 0
rect -56 -2 -5 0
rect -3 -2 6 0
rect 8 -2 46 0
rect 48 -2 56 0
rect 58 -2 87 0
rect 89 -2 140 0
rect 142 -2 151 0
rect 153 -2 161 0
rect 163 -2 192 0
rect 194 -2 245 0
rect 247 -2 256 0
rect 258 -2 296 0
rect 298 -2 306 0
rect 308 -2 337 0
rect 339 -2 390 0
rect 392 -2 401 0
rect 403 -2 411 0
rect 413 -2 442 0
rect 444 -2 495 0
rect 497 -2 506 0
rect 508 -2 546 0
rect 548 -2 556 0
rect 558 -2 587 0
rect 589 -2 640 0
rect 642 -2 651 0
rect 653 -2 661 0
rect 663 -2 692 0
rect 694 -2 745 0
rect 747 -2 753 0
rect -251 -3 753 -2
rect -207 -12 -195 -8
rect -207 -14 -205 -12
rect -203 -14 -195 -12
rect -130 -10 -106 -9
rect -247 -17 -242 -15
rect -247 -19 -245 -17
rect -243 -19 -242 -17
rect -247 -21 -242 -19
rect -247 -40 -243 -21
rect -215 -25 -211 -16
rect -207 -25 -203 -14
rect -130 -12 -128 -10
rect -126 -12 -106 -10
rect -130 -13 -106 -12
rect -247 -42 -245 -40
rect -247 -47 -243 -42
rect -247 -49 -245 -47
rect -232 -26 -203 -25
rect -232 -28 -228 -26
rect -226 -28 -203 -26
rect -232 -29 -203 -28
rect -232 -35 -218 -33
rect -216 -35 -211 -33
rect -232 -37 -211 -35
rect -215 -43 -211 -37
rect -215 -45 -214 -43
rect -212 -45 -211 -43
rect -215 -46 -211 -45
rect -207 -34 -203 -29
rect -183 -17 -178 -16
rect -183 -19 -182 -17
rect -180 -19 -178 -17
rect -183 -25 -178 -19
rect -207 -36 -202 -34
rect -207 -38 -205 -36
rect -203 -38 -202 -36
rect -207 -43 -202 -38
rect -207 -45 -205 -43
rect -203 -45 -202 -43
rect -192 -26 -178 -25
rect -192 -28 -188 -26
rect -186 -28 -178 -26
rect -192 -29 -178 -28
rect -158 -17 -145 -16
rect -158 -19 -155 -17
rect -153 -19 -145 -17
rect -158 -21 -145 -19
rect -110 -17 -106 -13
rect -158 -22 -148 -21
rect -150 -23 -148 -22
rect -146 -23 -145 -21
rect -166 -33 -161 -32
rect -184 -34 -171 -33
rect -167 -34 -161 -33
rect -184 -36 -178 -34
rect -176 -36 -164 -34
rect -162 -36 -161 -34
rect -184 -37 -161 -36
rect -175 -39 -161 -37
rect -150 -30 -145 -23
rect -110 -19 -109 -17
rect -107 -19 -106 -17
rect -207 -47 -202 -45
rect -247 -53 -234 -49
rect -247 -54 -243 -53
rect -175 -46 -171 -39
rect -166 -48 -161 -39
rect -166 -54 -154 -48
rect -110 -41 -106 -19
rect -122 -43 -106 -41
rect -122 -45 -120 -43
rect -118 -45 -106 -43
rect -122 -46 -106 -45
rect -102 -12 -90 -8
rect -102 -14 -100 -12
rect -98 -14 -90 -12
rect -25 -10 -1 -9
rect -102 -34 -98 -14
rect -25 -12 -23 -10
rect -21 -12 -1 -10
rect -25 -13 -1 -12
rect -78 -17 -73 -16
rect -78 -19 -77 -17
rect -75 -19 -73 -17
rect -78 -25 -73 -19
rect -102 -36 -97 -34
rect -102 -38 -100 -36
rect -98 -38 -97 -36
rect -102 -43 -97 -38
rect -102 -45 -100 -43
rect -98 -45 -97 -43
rect -87 -26 -73 -25
rect -87 -28 -83 -26
rect -81 -28 -73 -26
rect -87 -29 -73 -28
rect -53 -17 -40 -16
rect -53 -19 -50 -17
rect -48 -19 -40 -17
rect -53 -21 -40 -19
rect -53 -22 -43 -21
rect -45 -23 -43 -22
rect -41 -23 -40 -21
rect -61 -33 -56 -32
rect -79 -34 -66 -33
rect -62 -34 -56 -33
rect -79 -36 -73 -34
rect -71 -35 -59 -34
rect -71 -36 -67 -35
rect -79 -37 -67 -36
rect -65 -36 -59 -35
rect -57 -36 -56 -34
rect -65 -37 -56 -36
rect -70 -39 -56 -37
rect -45 -30 -40 -23
rect -102 -47 -97 -45
rect -70 -46 -66 -39
rect -61 -48 -56 -39
rect -61 -54 -49 -48
rect -5 -41 -1 -13
rect 43 -12 55 -8
rect 43 -14 45 -12
rect 47 -14 55 -12
rect 120 -10 144 -9
rect -17 -43 -1 -41
rect -17 -45 -15 -43
rect -13 -45 -1 -43
rect -17 -46 -1 -45
rect 3 -17 8 -15
rect 3 -19 5 -17
rect 7 -19 8 -17
rect 3 -21 8 -19
rect 3 -35 7 -21
rect 3 -37 4 -35
rect 6 -37 7 -35
rect 3 -40 7 -37
rect 35 -25 39 -16
rect 43 -25 47 -14
rect 120 -12 122 -10
rect 124 -12 144 -10
rect 120 -13 144 -12
rect 3 -42 5 -40
rect 3 -47 7 -42
rect 3 -49 5 -47
rect 18 -26 47 -25
rect 18 -28 22 -26
rect 24 -28 47 -26
rect 18 -29 47 -28
rect 18 -35 32 -33
rect 34 -35 39 -33
rect 18 -37 39 -35
rect 35 -43 39 -37
rect 35 -45 36 -43
rect 38 -45 39 -43
rect 35 -46 39 -45
rect 43 -34 47 -29
rect 67 -17 72 -16
rect 67 -19 68 -17
rect 70 -19 72 -17
rect 67 -25 72 -19
rect 43 -36 48 -34
rect 43 -38 45 -36
rect 47 -38 48 -36
rect 43 -43 48 -38
rect 43 -45 45 -43
rect 47 -45 48 -43
rect 58 -26 72 -25
rect 58 -28 62 -26
rect 64 -28 72 -26
rect 58 -29 72 -28
rect 92 -17 105 -16
rect 92 -19 95 -17
rect 97 -19 105 -17
rect 92 -21 105 -19
rect 140 -17 144 -13
rect 92 -22 102 -21
rect 100 -23 102 -22
rect 104 -23 105 -21
rect 84 -33 89 -32
rect 66 -34 79 -33
rect 83 -34 89 -33
rect 66 -36 72 -34
rect 74 -36 86 -34
rect 88 -36 89 -34
rect 66 -37 89 -36
rect 75 -39 89 -37
rect 100 -30 105 -23
rect 140 -19 141 -17
rect 143 -19 144 -17
rect 43 -47 48 -45
rect 3 -53 16 -49
rect 3 -54 7 -53
rect 75 -46 79 -39
rect 84 -48 89 -39
rect 84 -54 96 -48
rect 140 -41 144 -19
rect 128 -43 144 -41
rect 128 -45 130 -43
rect 132 -45 144 -43
rect 128 -46 144 -45
rect 148 -12 160 -8
rect 148 -14 150 -12
rect 152 -14 160 -12
rect 225 -10 249 -9
rect 148 -34 152 -14
rect 225 -12 227 -10
rect 229 -12 249 -10
rect 225 -13 249 -12
rect 172 -17 177 -16
rect 172 -19 173 -17
rect 175 -19 177 -17
rect 172 -25 177 -19
rect 148 -36 153 -34
rect 148 -38 150 -36
rect 152 -38 153 -36
rect 148 -43 153 -38
rect 148 -45 150 -43
rect 152 -45 153 -43
rect 163 -26 177 -25
rect 163 -28 167 -26
rect 169 -28 177 -26
rect 163 -29 177 -28
rect 197 -17 210 -16
rect 197 -19 200 -17
rect 202 -19 210 -17
rect 197 -21 210 -19
rect 197 -22 207 -21
rect 205 -23 207 -22
rect 209 -23 210 -21
rect 189 -33 194 -32
rect 171 -34 184 -33
rect 188 -34 194 -33
rect 171 -36 177 -34
rect 179 -35 191 -34
rect 179 -36 185 -35
rect 171 -37 185 -36
rect 187 -36 191 -35
rect 193 -36 194 -34
rect 187 -37 194 -36
rect 180 -39 194 -37
rect 205 -30 210 -23
rect 148 -47 153 -45
rect 180 -46 184 -39
rect 189 -48 194 -39
rect 189 -54 201 -48
rect 245 -41 249 -13
rect 293 -12 305 -8
rect 293 -14 295 -12
rect 297 -14 305 -12
rect 370 -10 394 -9
rect 233 -43 249 -41
rect 233 -45 235 -43
rect 237 -45 249 -43
rect 233 -46 249 -45
rect 253 -17 258 -15
rect 253 -19 255 -17
rect 257 -19 258 -17
rect 253 -21 258 -19
rect 253 -35 257 -21
rect 253 -37 254 -35
rect 256 -37 257 -35
rect 253 -40 257 -37
rect 285 -25 289 -16
rect 293 -25 297 -14
rect 370 -12 372 -10
rect 374 -12 394 -10
rect 370 -13 394 -12
rect 253 -42 255 -40
rect 253 -47 257 -42
rect 253 -49 255 -47
rect 268 -26 297 -25
rect 268 -28 272 -26
rect 274 -28 297 -26
rect 268 -29 297 -28
rect 268 -35 282 -33
rect 284 -35 289 -33
rect 268 -37 289 -35
rect 285 -43 289 -37
rect 285 -45 286 -43
rect 288 -45 289 -43
rect 285 -46 289 -45
rect 293 -34 297 -29
rect 317 -17 322 -16
rect 317 -19 318 -17
rect 320 -19 322 -17
rect 317 -25 322 -19
rect 293 -36 298 -34
rect 293 -38 295 -36
rect 297 -38 298 -36
rect 293 -43 298 -38
rect 293 -45 295 -43
rect 297 -45 298 -43
rect 308 -26 322 -25
rect 308 -28 312 -26
rect 314 -28 322 -26
rect 308 -29 322 -28
rect 342 -17 355 -16
rect 342 -19 345 -17
rect 347 -19 355 -17
rect 342 -21 355 -19
rect 390 -17 394 -13
rect 342 -22 352 -21
rect 350 -23 352 -22
rect 354 -23 355 -21
rect 334 -33 339 -32
rect 316 -34 329 -33
rect 333 -34 339 -33
rect 316 -36 322 -34
rect 324 -36 336 -34
rect 338 -36 339 -34
rect 316 -37 339 -36
rect 325 -39 339 -37
rect 350 -30 355 -23
rect 390 -19 391 -17
rect 393 -19 394 -17
rect 293 -47 298 -45
rect 253 -53 266 -49
rect 253 -54 257 -53
rect 325 -46 329 -39
rect 334 -48 339 -39
rect 334 -54 346 -48
rect 390 -41 394 -19
rect 378 -43 394 -41
rect 378 -45 380 -43
rect 382 -45 394 -43
rect 378 -46 394 -45
rect 398 -12 410 -8
rect 398 -14 400 -12
rect 402 -14 410 -12
rect 475 -10 499 -9
rect 398 -34 402 -14
rect 475 -12 477 -10
rect 479 -12 499 -10
rect 475 -13 499 -12
rect 422 -17 427 -16
rect 422 -19 423 -17
rect 425 -19 427 -17
rect 422 -25 427 -19
rect 398 -36 403 -34
rect 398 -38 400 -36
rect 402 -38 403 -36
rect 398 -43 403 -38
rect 398 -45 400 -43
rect 402 -45 403 -43
rect 413 -26 427 -25
rect 413 -28 417 -26
rect 419 -28 427 -26
rect 413 -29 427 -28
rect 447 -17 460 -16
rect 447 -19 450 -17
rect 452 -19 460 -17
rect 447 -21 460 -19
rect 447 -22 457 -21
rect 455 -23 457 -22
rect 459 -23 460 -21
rect 439 -33 444 -32
rect 421 -34 434 -33
rect 438 -34 444 -33
rect 421 -36 427 -34
rect 429 -35 441 -34
rect 429 -36 435 -35
rect 421 -37 435 -36
rect 437 -36 441 -35
rect 443 -36 444 -34
rect 437 -37 444 -36
rect 430 -39 444 -37
rect 455 -30 460 -23
rect 398 -47 403 -45
rect 430 -46 434 -39
rect 439 -48 444 -39
rect 439 -54 451 -48
rect 495 -41 499 -13
rect 543 -12 555 -8
rect 543 -14 545 -12
rect 547 -14 555 -12
rect 620 -10 644 -9
rect 483 -43 499 -41
rect 483 -45 485 -43
rect 487 -45 499 -43
rect 483 -46 499 -45
rect 503 -17 508 -15
rect 503 -19 505 -17
rect 507 -19 508 -17
rect 503 -21 508 -19
rect 503 -35 507 -21
rect 503 -37 504 -35
rect 506 -37 507 -35
rect 503 -40 507 -37
rect 535 -25 539 -16
rect 543 -25 547 -14
rect 620 -12 622 -10
rect 624 -12 644 -10
rect 620 -13 644 -12
rect 503 -42 505 -40
rect 503 -47 507 -42
rect 503 -49 505 -47
rect 518 -26 547 -25
rect 518 -28 522 -26
rect 524 -28 547 -26
rect 518 -29 547 -28
rect 518 -35 532 -33
rect 534 -35 539 -33
rect 518 -37 539 -35
rect 535 -43 539 -37
rect 535 -45 536 -43
rect 538 -45 539 -43
rect 535 -46 539 -45
rect 543 -34 547 -29
rect 567 -17 572 -16
rect 567 -19 568 -17
rect 570 -19 572 -17
rect 567 -25 572 -19
rect 543 -36 548 -34
rect 543 -38 545 -36
rect 547 -38 548 -36
rect 543 -43 548 -38
rect 543 -45 545 -43
rect 547 -45 548 -43
rect 558 -26 572 -25
rect 558 -28 562 -26
rect 564 -28 572 -26
rect 558 -29 572 -28
rect 592 -17 605 -16
rect 592 -19 595 -17
rect 597 -19 605 -17
rect 592 -21 605 -19
rect 640 -17 644 -13
rect 592 -22 602 -21
rect 600 -23 602 -22
rect 604 -23 605 -21
rect 584 -33 589 -32
rect 566 -34 579 -33
rect 583 -34 589 -33
rect 566 -36 572 -34
rect 574 -36 586 -34
rect 588 -36 589 -34
rect 566 -37 589 -36
rect 575 -39 589 -37
rect 600 -30 605 -23
rect 640 -19 641 -17
rect 643 -19 644 -17
rect 543 -47 548 -45
rect 503 -53 516 -49
rect 503 -54 507 -53
rect 575 -46 579 -39
rect 584 -48 589 -39
rect 584 -54 596 -48
rect 640 -41 644 -19
rect 628 -43 644 -41
rect 628 -45 630 -43
rect 632 -45 644 -43
rect 628 -46 644 -45
rect 648 -12 660 -8
rect 648 -14 650 -12
rect 652 -14 660 -12
rect 725 -10 749 -9
rect 648 -34 652 -14
rect 725 -12 727 -10
rect 729 -12 749 -10
rect 725 -13 749 -12
rect 672 -17 677 -16
rect 672 -19 673 -17
rect 675 -19 677 -17
rect 672 -25 677 -19
rect 648 -36 653 -34
rect 648 -38 650 -36
rect 652 -38 653 -36
rect 648 -43 653 -38
rect 648 -45 650 -43
rect 652 -45 653 -43
rect 663 -26 677 -25
rect 663 -28 667 -26
rect 669 -28 677 -26
rect 663 -29 677 -28
rect 697 -17 710 -16
rect 697 -19 700 -17
rect 702 -19 710 -17
rect 697 -21 710 -19
rect 697 -22 707 -21
rect 705 -23 707 -22
rect 709 -23 710 -21
rect 689 -33 694 -32
rect 671 -34 684 -33
rect 688 -34 694 -33
rect 671 -36 677 -34
rect 679 -36 691 -34
rect 693 -36 694 -34
rect 671 -37 694 -36
rect 680 -39 694 -37
rect 705 -30 710 -23
rect 648 -47 653 -45
rect 680 -46 684 -39
rect 689 -48 694 -39
rect 689 -54 701 -48
rect 745 -41 749 -13
rect 733 -43 749 -41
rect 733 -45 735 -43
rect 737 -45 749 -43
rect 733 -46 749 -45
rect -251 -60 753 -59
rect -251 -62 -244 -60
rect -242 -62 -204 -60
rect -202 -62 -130 -60
rect -128 -62 -99 -60
rect -97 -62 -25 -60
rect -23 -62 6 -60
rect 8 -62 46 -60
rect 48 -62 120 -60
rect 122 -62 151 -60
rect 153 -62 225 -60
rect 227 -62 256 -60
rect 258 -62 296 -60
rect 298 -62 370 -60
rect 372 -62 401 -60
rect 403 -62 475 -60
rect 477 -62 506 -60
rect 508 -62 546 -60
rect 548 -62 620 -60
rect 622 -62 651 -60
rect 653 -62 725 -60
rect 727 -62 753 -60
rect -251 -67 753 -62
<< alu2 >>
rect 51 127 183 128
rect 51 125 52 127
rect 54 125 153 127
rect 155 125 180 127
rect 182 125 183 127
rect 51 124 183 125
rect 256 127 388 128
rect 256 125 257 127
rect 259 125 358 127
rect 360 125 385 127
rect 387 125 388 127
rect 256 124 388 125
rect 34 118 40 119
rect 34 116 37 118
rect 39 116 40 118
rect 11 102 23 103
rect 11 100 20 102
rect 22 100 23 102
rect 11 98 23 100
rect 11 25 16 98
rect 34 38 40 116
rect 76 118 80 119
rect 76 116 77 118
rect 79 116 80 118
rect 59 103 63 104
rect 59 101 60 103
rect 62 101 63 103
rect 59 77 63 101
rect 51 73 63 77
rect 51 55 55 73
rect 51 53 52 55
rect 54 53 55 55
rect 51 52 55 53
rect 34 36 35 38
rect 37 36 40 38
rect 34 35 40 36
rect 59 46 63 47
rect 59 44 60 46
rect 62 44 63 46
rect 59 25 63 44
rect 76 38 80 116
rect 203 115 207 119
rect 203 113 204 115
rect 206 113 207 115
rect 90 104 175 105
rect 90 102 91 104
rect 93 102 172 104
rect 174 102 175 104
rect 90 101 175 102
rect 203 78 207 113
rect 239 118 245 119
rect 239 116 242 118
rect 244 116 245 118
rect 147 73 207 78
rect 216 102 228 103
rect 216 100 225 102
rect 227 100 228 102
rect 216 98 228 100
rect 147 62 152 73
rect 147 60 148 62
rect 150 60 152 62
rect 147 58 152 60
rect 76 36 77 38
rect 79 36 80 38
rect 76 35 80 36
rect 91 29 156 30
rect 91 27 92 29
rect 94 27 124 29
rect 126 27 151 29
rect 153 27 156 29
rect 91 26 156 27
rect 91 25 129 26
rect 216 25 221 98
rect 239 38 245 116
rect 281 118 285 119
rect 281 116 282 118
rect 284 116 285 118
rect 264 103 268 104
rect 264 101 265 103
rect 267 101 268 103
rect 264 77 268 101
rect 256 73 268 77
rect 256 55 260 73
rect 256 53 257 55
rect 259 53 260 55
rect 256 52 260 53
rect 239 36 240 38
rect 242 36 245 38
rect 239 35 245 36
rect 264 46 268 47
rect 264 44 265 46
rect 267 44 268 46
rect 264 25 268 44
rect 281 38 285 116
rect 408 115 412 119
rect 408 113 409 115
rect 411 113 412 115
rect 295 104 380 105
rect 295 102 296 104
rect 298 102 377 104
rect 379 102 380 104
rect 295 101 380 102
rect 408 78 412 113
rect 352 73 412 78
rect 352 62 357 73
rect 352 60 353 62
rect 355 60 357 62
rect 352 58 357 60
rect 281 36 282 38
rect 284 36 285 38
rect 281 35 285 36
rect 296 29 361 30
rect 296 27 297 29
rect 299 27 329 29
rect 331 27 356 29
rect 358 27 361 29
rect 296 26 361 27
rect 296 25 334 26
rect 11 21 63 25
rect 216 21 268 25
rect -183 -17 -150 -16
rect -183 -19 -182 -17
rect -180 -19 -155 -17
rect -153 -19 -150 -17
rect -183 -20 -150 -19
rect -110 -17 -45 -16
rect -110 -19 -109 -17
rect -107 -19 -77 -17
rect -75 -19 -50 -17
rect -48 -19 -45 -17
rect -110 -20 -45 -19
rect 67 -17 100 -16
rect 67 -19 68 -17
rect 70 -19 95 -17
rect 97 -19 100 -17
rect 67 -20 100 -19
rect 140 -17 205 -16
rect 140 -19 141 -17
rect 143 -19 173 -17
rect 175 -19 200 -17
rect 202 -19 205 -17
rect 140 -20 205 -19
rect 317 -17 350 -16
rect 317 -19 318 -17
rect 320 -19 345 -17
rect 347 -19 350 -17
rect 317 -20 350 -19
rect 390 -17 455 -16
rect 390 -19 391 -17
rect 393 -19 423 -17
rect 425 -19 450 -17
rect 452 -19 455 -17
rect 390 -20 455 -19
rect 567 -17 600 -16
rect 567 -19 568 -17
rect 570 -19 595 -17
rect 597 -19 600 -17
rect 567 -20 600 -19
rect 640 -17 705 -16
rect 640 -19 641 -17
rect 643 -19 673 -17
rect 675 -19 700 -17
rect 702 -19 705 -17
rect 640 -20 705 -19
rect -68 -35 7 -34
rect -68 -37 -67 -35
rect -65 -37 4 -35
rect 6 -37 7 -35
rect -68 -38 7 -37
rect 184 -35 257 -34
rect 184 -37 185 -35
rect 187 -37 254 -35
rect 256 -37 257 -35
rect 184 -38 257 -37
rect 434 -35 507 -34
rect 434 -37 435 -35
rect 437 -37 504 -35
rect 506 -37 507 -35
rect 434 -38 507 -37
rect -215 -43 -97 -42
rect -215 -45 -214 -43
rect -212 -45 -100 -43
rect -98 -45 -97 -43
rect -215 -46 -97 -45
rect 35 -43 153 -42
rect 35 -45 36 -43
rect 38 -45 150 -43
rect 152 -45 153 -43
rect 35 -46 153 -45
rect 285 -43 403 -42
rect 285 -45 286 -43
rect 288 -45 400 -43
rect 402 -45 403 -43
rect 285 -46 403 -45
rect 535 -43 653 -42
rect 535 -45 536 -43
rect 538 -45 650 -43
rect 652 -45 653 -43
rect 535 -46 653 -45
<< ptie >>
rect 48 144 54 146
rect 48 142 50 144
rect 52 142 54 144
rect 48 140 54 142
rect 88 144 94 146
rect 88 142 90 144
rect 92 142 94 144
rect 88 140 94 142
rect 159 144 165 146
rect 159 142 161 144
rect 163 142 165 144
rect 159 140 165 142
rect 200 144 206 146
rect 200 142 202 144
rect 204 142 206 144
rect 200 140 206 142
rect 253 144 259 146
rect 253 142 255 144
rect 257 142 259 144
rect 253 140 259 142
rect 293 144 299 146
rect 293 142 295 144
rect 297 142 299 144
rect 293 140 299 142
rect 364 144 370 146
rect 364 142 366 144
rect 368 142 370 144
rect 364 140 370 142
rect 405 144 411 146
rect 405 142 407 144
rect 409 142 411 144
rect 405 140 411 142
rect 20 12 26 14
rect 20 10 22 12
rect 24 10 26 12
rect 20 8 26 10
rect 88 12 94 14
rect 88 10 90 12
rect 92 10 94 12
rect 88 8 94 10
rect 100 12 106 14
rect 100 10 102 12
rect 104 10 106 12
rect 100 8 106 10
rect 141 12 147 14
rect 141 10 143 12
rect 145 10 147 12
rect 141 8 147 10
rect 225 12 231 14
rect 225 10 227 12
rect 229 10 231 12
rect 225 8 231 10
rect 293 12 299 14
rect 293 10 295 12
rect 297 10 299 12
rect 293 8 299 10
rect 305 12 311 14
rect 305 10 307 12
rect 309 10 311 12
rect 305 8 311 10
rect 346 12 352 14
rect 346 10 348 12
rect 350 10 352 12
rect 346 8 352 10
rect -246 0 -240 2
rect -246 -2 -244 0
rect -242 -2 -240 0
rect -206 0 -200 2
rect -206 -2 -204 0
rect -202 -2 -200 0
rect -246 -4 -240 -2
rect -206 -4 -200 -2
rect -165 0 -159 2
rect -165 -2 -163 0
rect -161 -2 -159 0
rect -165 -4 -159 -2
rect -101 0 -95 2
rect -101 -2 -99 0
rect -97 -2 -95 0
rect -101 -4 -95 -2
rect -60 0 -54 2
rect -60 -2 -58 0
rect -56 -2 -54 0
rect -60 -4 -54 -2
rect 4 0 10 2
rect 4 -2 6 0
rect 8 -2 10 0
rect 44 0 50 2
rect 44 -2 46 0
rect 48 -2 50 0
rect 4 -4 10 -2
rect 44 -4 50 -2
rect 85 0 91 2
rect 85 -2 87 0
rect 89 -2 91 0
rect 85 -4 91 -2
rect 149 0 155 2
rect 149 -2 151 0
rect 153 -2 155 0
rect 149 -4 155 -2
rect 190 0 196 2
rect 190 -2 192 0
rect 194 -2 196 0
rect 190 -4 196 -2
rect 254 0 260 2
rect 254 -2 256 0
rect 258 -2 260 0
rect 294 0 300 2
rect 294 -2 296 0
rect 298 -2 300 0
rect 254 -4 260 -2
rect 294 -4 300 -2
rect 335 0 341 2
rect 335 -2 337 0
rect 339 -2 341 0
rect 335 -4 341 -2
rect 399 0 405 2
rect 399 -2 401 0
rect 403 -2 405 0
rect 399 -4 405 -2
rect 440 0 446 2
rect 440 -2 442 0
rect 444 -2 446 0
rect 440 -4 446 -2
rect 504 0 510 2
rect 504 -2 506 0
rect 508 -2 510 0
rect 544 0 550 2
rect 544 -2 546 0
rect 548 -2 550 0
rect 504 -4 510 -2
rect 544 -4 550 -2
rect 585 0 591 2
rect 585 -2 587 0
rect 589 -2 591 0
rect 585 -4 591 -2
rect 649 0 655 2
rect 649 -2 651 0
rect 653 -2 655 0
rect 649 -4 655 -2
rect 690 0 696 2
rect 690 -2 692 0
rect 694 -2 696 0
rect 690 -4 696 -2
<< ntie >>
rect 48 84 54 86
rect 48 82 50 84
rect 52 82 54 84
rect 48 80 54 82
rect 88 84 94 86
rect 88 82 90 84
rect 92 82 94 84
rect 126 84 132 86
rect 88 80 94 82
rect 126 82 128 84
rect 130 82 132 84
rect 200 84 206 86
rect 126 80 132 82
rect 200 82 202 84
rect 204 82 206 84
rect 200 80 206 82
rect 253 84 259 86
rect 253 82 255 84
rect 257 82 259 84
rect 253 80 259 82
rect 293 84 299 86
rect 293 82 295 84
rect 297 82 299 84
rect 331 84 337 86
rect 293 80 299 82
rect 331 82 333 84
rect 335 82 337 84
rect 405 84 411 86
rect 331 80 337 82
rect 405 82 407 84
rect 409 82 411 84
rect 405 80 411 82
rect 20 72 26 74
rect 20 70 22 72
rect 24 70 26 72
rect 20 68 26 70
rect 88 72 94 74
rect 88 70 90 72
rect 92 70 94 72
rect 88 68 94 70
rect 100 72 106 74
rect 100 70 102 72
rect 104 70 106 72
rect 174 72 180 74
rect 100 68 106 70
rect 174 70 176 72
rect 178 70 180 72
rect 225 72 231 74
rect 174 68 180 70
rect 225 70 227 72
rect 229 70 231 72
rect 225 68 231 70
rect 293 72 299 74
rect 293 70 295 72
rect 297 70 299 72
rect 293 68 299 70
rect 305 72 311 74
rect 305 70 307 72
rect 309 70 311 72
rect 379 72 385 74
rect 305 68 311 70
rect 379 70 381 72
rect 383 70 385 72
rect 379 68 385 70
rect -246 -60 -240 -58
rect -246 -62 -244 -60
rect -242 -62 -240 -60
rect -206 -60 -200 -58
rect -246 -64 -240 -62
rect -206 -62 -204 -60
rect -202 -62 -200 -60
rect -132 -60 -126 -58
rect -206 -64 -200 -62
rect -132 -62 -130 -60
rect -128 -62 -126 -60
rect -101 -60 -95 -58
rect -132 -64 -126 -62
rect -101 -62 -99 -60
rect -97 -62 -95 -60
rect -27 -60 -21 -58
rect -101 -64 -95 -62
rect -27 -62 -25 -60
rect -23 -62 -21 -60
rect 4 -60 10 -58
rect -27 -64 -21 -62
rect 4 -62 6 -60
rect 8 -62 10 -60
rect 44 -60 50 -58
rect 4 -64 10 -62
rect 44 -62 46 -60
rect 48 -62 50 -60
rect 118 -60 124 -58
rect 44 -64 50 -62
rect 118 -62 120 -60
rect 122 -62 124 -60
rect 149 -60 155 -58
rect 118 -64 124 -62
rect 149 -62 151 -60
rect 153 -62 155 -60
rect 223 -60 229 -58
rect 149 -64 155 -62
rect 223 -62 225 -60
rect 227 -62 229 -60
rect 254 -60 260 -58
rect 223 -64 229 -62
rect 254 -62 256 -60
rect 258 -62 260 -60
rect 294 -60 300 -58
rect 254 -64 260 -62
rect 294 -62 296 -60
rect 298 -62 300 -60
rect 368 -60 374 -58
rect 294 -64 300 -62
rect 368 -62 370 -60
rect 372 -62 374 -60
rect 399 -60 405 -58
rect 368 -64 374 -62
rect 399 -62 401 -60
rect 403 -62 405 -60
rect 473 -60 479 -58
rect 399 -64 405 -62
rect 473 -62 475 -60
rect 477 -62 479 -60
rect 504 -60 510 -58
rect 473 -64 479 -62
rect 504 -62 506 -60
rect 508 -62 510 -60
rect 544 -60 550 -58
rect 504 -64 510 -62
rect 544 -62 546 -60
rect 548 -62 550 -60
rect 618 -60 624 -58
rect 544 -64 550 -62
rect 618 -62 620 -60
rect 622 -62 624 -60
rect 649 -60 655 -58
rect 618 -64 624 -62
rect 649 -62 651 -60
rect 653 -62 655 -60
rect 723 -60 729 -58
rect 649 -64 655 -62
rect 723 -62 725 -60
rect 727 -62 729 -60
rect 723 -64 729 -62
<< nmos >>
rect 26 125 28 136
rect 33 125 35 136
rect 46 125 48 134
rect 66 125 68 136
rect 73 125 75 136
rect 86 125 88 134
rect 114 128 116 140
rect 121 128 123 140
rect 131 128 133 137
rect 141 128 143 137
rect 157 123 159 132
rect 178 125 180 136
rect 185 125 187 136
rect 198 125 200 134
rect 231 125 233 136
rect 238 125 240 136
rect 251 125 253 134
rect 271 125 273 136
rect 278 125 280 136
rect 291 125 293 134
rect 319 128 321 140
rect 326 128 328 140
rect 336 128 338 137
rect 346 128 348 137
rect 362 123 364 132
rect 383 125 385 136
rect 390 125 392 136
rect 403 125 405 134
rect 26 20 28 29
rect 39 18 41 29
rect 46 18 48 29
rect 66 18 68 29
rect 73 18 75 29
rect 86 20 88 29
rect 106 20 108 29
rect 119 18 121 29
rect 126 18 128 29
rect 147 22 149 31
rect 163 17 165 26
rect 173 17 175 26
rect 183 14 185 26
rect 190 14 192 26
rect 231 20 233 29
rect 244 18 246 29
rect 251 18 253 29
rect 271 18 273 29
rect 278 18 280 29
rect 291 20 293 29
rect 311 20 313 29
rect 324 18 326 29
rect 331 18 333 29
rect 352 22 354 31
rect 368 17 370 26
rect 378 17 380 26
rect 388 14 390 26
rect 395 14 397 26
rect -240 -21 -238 -12
rect -230 -21 -228 -15
rect -220 -21 -218 -15
rect -200 -19 -198 -10
rect -187 -19 -185 -8
rect -180 -19 -178 -8
rect -159 -21 -157 -12
rect -143 -16 -141 -7
rect -133 -16 -131 -7
rect -123 -16 -121 -4
rect -116 -16 -114 -4
rect -95 -19 -93 -10
rect -82 -19 -80 -8
rect -75 -19 -73 -8
rect -54 -21 -52 -12
rect -38 -16 -36 -7
rect -28 -16 -26 -7
rect -18 -16 -16 -4
rect -11 -16 -9 -4
rect 10 -21 12 -12
rect 20 -21 22 -15
rect 30 -21 32 -15
rect 50 -19 52 -10
rect 63 -19 65 -8
rect 70 -19 72 -8
rect 91 -21 93 -12
rect 107 -16 109 -7
rect 117 -16 119 -7
rect 127 -16 129 -4
rect 134 -16 136 -4
rect 155 -19 157 -10
rect 168 -19 170 -8
rect 175 -19 177 -8
rect 196 -21 198 -12
rect 212 -16 214 -7
rect 222 -16 224 -7
rect 232 -16 234 -4
rect 239 -16 241 -4
rect 260 -21 262 -12
rect 270 -21 272 -15
rect 280 -21 282 -15
rect 300 -19 302 -10
rect 313 -19 315 -8
rect 320 -19 322 -8
rect 341 -21 343 -12
rect 357 -16 359 -7
rect 367 -16 369 -7
rect 377 -16 379 -4
rect 384 -16 386 -4
rect 405 -19 407 -10
rect 418 -19 420 -8
rect 425 -19 427 -8
rect 446 -21 448 -12
rect 462 -16 464 -7
rect 472 -16 474 -7
rect 482 -16 484 -4
rect 489 -16 491 -4
rect 510 -21 512 -12
rect 520 -21 522 -15
rect 530 -21 532 -15
rect 550 -19 552 -10
rect 563 -19 565 -8
rect 570 -19 572 -8
rect 591 -21 593 -12
rect 607 -16 609 -7
rect 617 -16 619 -7
rect 627 -16 629 -4
rect 634 -16 636 -4
rect 655 -19 657 -10
rect 668 -19 670 -8
rect 675 -19 677 -8
rect 696 -21 698 -12
rect 712 -16 714 -7
rect 722 -16 724 -7
rect 732 -16 734 -4
rect 739 -16 741 -4
<< pmos >>
rect 26 90 28 103
rect 36 90 38 103
rect 46 92 48 110
rect 66 90 68 103
rect 76 90 78 103
rect 86 92 88 110
rect 113 83 115 110
rect 123 92 125 110
rect 133 92 135 110
rect 149 83 151 110
rect 178 90 180 103
rect 188 90 190 103
rect 198 92 200 110
rect 231 90 233 103
rect 241 90 243 103
rect 251 92 253 110
rect 271 90 273 103
rect 281 90 283 103
rect 291 92 293 110
rect 318 83 320 110
rect 328 92 330 110
rect 338 92 340 110
rect 354 83 356 110
rect 383 90 385 103
rect 393 90 395 103
rect 403 92 405 110
rect 26 44 28 62
rect 36 51 38 64
rect 46 51 48 64
rect 66 51 68 64
rect 76 51 78 64
rect 86 44 88 62
rect 106 44 108 62
rect 116 51 118 64
rect 126 51 128 64
rect 155 44 157 71
rect 171 44 173 62
rect 181 44 183 62
rect 191 44 193 71
rect 231 44 233 62
rect 241 51 243 64
rect 251 51 253 64
rect 271 51 273 64
rect 281 51 283 64
rect 291 44 293 62
rect 311 44 313 62
rect 321 51 323 64
rect 331 51 333 64
rect 360 44 362 71
rect 376 44 378 62
rect 386 44 388 62
rect 396 44 398 71
rect -240 -51 -238 -33
rect -227 -61 -225 -40
rect -220 -61 -218 -40
rect -200 -52 -198 -34
rect -190 -54 -188 -41
rect -180 -54 -178 -41
rect -151 -61 -149 -34
rect -135 -52 -133 -34
rect -125 -52 -123 -34
rect -115 -61 -113 -34
rect -95 -52 -93 -34
rect -85 -54 -83 -41
rect -75 -54 -73 -41
rect -46 -61 -44 -34
rect -30 -52 -28 -34
rect -20 -52 -18 -34
rect -10 -61 -8 -34
rect 10 -51 12 -33
rect 23 -61 25 -40
rect 30 -61 32 -40
rect 50 -52 52 -34
rect 60 -54 62 -41
rect 70 -54 72 -41
rect 99 -61 101 -34
rect 115 -52 117 -34
rect 125 -52 127 -34
rect 135 -61 137 -34
rect 155 -52 157 -34
rect 165 -54 167 -41
rect 175 -54 177 -41
rect 204 -61 206 -34
rect 220 -52 222 -34
rect 230 -52 232 -34
rect 240 -61 242 -34
rect 260 -51 262 -33
rect 273 -61 275 -40
rect 280 -61 282 -40
rect 300 -52 302 -34
rect 310 -54 312 -41
rect 320 -54 322 -41
rect 349 -61 351 -34
rect 365 -52 367 -34
rect 375 -52 377 -34
rect 385 -61 387 -34
rect 405 -52 407 -34
rect 415 -54 417 -41
rect 425 -54 427 -41
rect 454 -61 456 -34
rect 470 -52 472 -34
rect 480 -52 482 -34
rect 490 -61 492 -34
rect 510 -51 512 -33
rect 523 -61 525 -40
rect 530 -61 532 -40
rect 550 -52 552 -34
rect 560 -54 562 -41
rect 570 -54 572 -41
rect 599 -61 601 -34
rect 615 -52 617 -34
rect 625 -52 627 -34
rect 635 -61 637 -34
rect 655 -52 657 -34
rect 665 -54 667 -41
rect 675 -54 677 -41
rect 704 -61 706 -34
rect 720 -52 722 -34
rect 730 -52 732 -34
rect 740 -61 742 -34
<< polyct0 >>
rect 44 116 46 118
rect 84 116 86 118
rect 115 115 117 117
rect 125 116 127 118
rect 196 116 198 118
rect 249 116 251 118
rect 289 116 291 118
rect 320 115 322 117
rect 330 116 332 118
rect 401 116 403 118
rect 28 36 30 38
rect 84 36 86 38
rect 108 36 110 38
rect 179 36 181 38
rect 189 37 191 39
rect 233 36 235 38
rect 289 36 291 38
rect 313 36 315 38
rect 384 36 386 38
rect 394 37 396 39
rect -238 -28 -236 -26
rect -198 -28 -196 -26
rect -127 -28 -125 -26
rect -117 -29 -115 -27
rect -93 -28 -91 -26
rect -22 -28 -20 -26
rect -12 -29 -10 -27
rect 12 -28 14 -26
rect 52 -28 54 -26
rect 123 -28 125 -26
rect 133 -29 135 -27
rect 157 -28 159 -26
rect 228 -28 230 -26
rect 238 -29 240 -27
rect 262 -28 264 -26
rect 302 -28 304 -26
rect 373 -28 375 -26
rect 383 -29 385 -27
rect 407 -28 409 -26
rect 478 -28 480 -26
rect 488 -29 490 -27
rect 512 -28 514 -26
rect 552 -28 554 -26
rect 623 -28 625 -26
rect 633 -29 635 -27
rect 657 -28 659 -26
rect 728 -28 730 -26
rect 738 -29 740 -27
<< polyct1 >>
rect 34 116 36 118
rect 24 108 26 110
rect 74 116 76 118
rect 146 121 148 123
rect 64 108 66 110
rect 186 116 188 118
rect 162 108 164 110
rect 176 108 178 110
rect 239 116 241 118
rect 229 108 231 110
rect 279 116 281 118
rect 351 121 353 123
rect 269 108 271 110
rect 391 116 393 118
rect 367 108 369 110
rect 381 108 383 110
rect 48 44 50 46
rect 64 44 66 46
rect 38 36 40 38
rect 74 36 76 38
rect 128 44 130 46
rect 142 44 144 46
rect 118 36 120 38
rect 253 44 255 46
rect 269 44 271 46
rect 158 31 160 33
rect 243 36 245 38
rect 279 36 281 38
rect 333 44 335 46
rect 347 44 349 46
rect 323 36 325 38
rect 363 31 365 33
rect -228 -28 -226 -26
rect -188 -28 -186 -26
rect -218 -35 -216 -33
rect -148 -23 -146 -21
rect -178 -36 -176 -34
rect -83 -28 -81 -26
rect -164 -36 -162 -34
rect -43 -23 -41 -21
rect -73 -36 -71 -34
rect 22 -28 24 -26
rect -59 -36 -57 -34
rect 62 -28 64 -26
rect 32 -35 34 -33
rect 102 -23 104 -21
rect 72 -36 74 -34
rect 167 -28 169 -26
rect 86 -36 88 -34
rect 207 -23 209 -21
rect 177 -36 179 -34
rect 272 -28 274 -26
rect 191 -36 193 -34
rect 312 -28 314 -26
rect 282 -35 284 -33
rect 352 -23 354 -21
rect 322 -36 324 -34
rect 417 -28 419 -26
rect 336 -36 338 -34
rect 457 -23 459 -21
rect 427 -36 429 -34
rect 522 -28 524 -26
rect 441 -36 443 -34
rect 562 -28 564 -26
rect 532 -35 534 -33
rect 602 -23 604 -21
rect 572 -36 574 -34
rect 667 -28 669 -26
rect 586 -36 588 -34
rect 707 -23 709 -21
rect 677 -36 679 -34
rect 691 -36 693 -34
<< ndifct0 >>
rect 21 132 23 134
rect 61 132 63 134
rect 136 130 138 132
rect 148 133 150 135
rect 173 132 175 134
rect 162 125 164 127
rect 226 132 228 134
rect 266 132 268 134
rect 341 130 343 132
rect 353 133 355 135
rect 378 132 380 134
rect 367 125 369 127
rect 51 20 53 22
rect 61 20 63 22
rect 142 27 144 29
rect 131 20 133 22
rect 156 19 158 21
rect 168 22 170 24
rect 256 20 258 22
rect 266 20 268 22
rect 347 27 349 29
rect 336 20 338 22
rect 361 19 363 21
rect 373 22 375 24
rect -234 -6 -232 -4
rect -215 -6 -213 -4
rect -225 -19 -223 -17
rect -175 -12 -173 -10
rect -150 -11 -148 -9
rect -164 -19 -162 -17
rect -138 -14 -136 -12
rect -70 -12 -68 -10
rect -45 -11 -43 -9
rect -59 -19 -57 -17
rect -33 -14 -31 -12
rect 16 -6 18 -4
rect 35 -6 37 -4
rect 25 -19 27 -17
rect 75 -12 77 -10
rect 100 -11 102 -9
rect 86 -19 88 -17
rect 112 -14 114 -12
rect 180 -12 182 -10
rect 205 -11 207 -9
rect 191 -19 193 -17
rect 217 -14 219 -12
rect 266 -6 268 -4
rect 285 -6 287 -4
rect 275 -19 277 -17
rect 325 -12 327 -10
rect 350 -11 352 -9
rect 336 -19 338 -17
rect 362 -14 364 -12
rect 430 -12 432 -10
rect 455 -11 457 -9
rect 441 -19 443 -17
rect 467 -14 469 -12
rect 516 -6 518 -4
rect 535 -6 537 -4
rect 525 -19 527 -17
rect 575 -12 577 -10
rect 600 -11 602 -9
rect 586 -19 588 -17
rect 612 -14 614 -12
rect 680 -12 682 -10
rect 705 -11 707 -9
rect 691 -19 693 -17
rect 717 -14 719 -12
<< ndifct1 >>
rect 40 142 42 144
rect 80 142 82 144
rect 108 142 110 144
rect 51 130 53 132
rect 91 130 93 132
rect 192 142 194 144
rect 126 132 128 134
rect 245 142 247 144
rect 285 142 287 144
rect 203 130 205 132
rect 313 142 315 144
rect 256 130 258 132
rect 296 130 298 132
rect 397 142 399 144
rect 331 132 333 134
rect 408 130 410 132
rect 21 22 23 24
rect 91 22 93 24
rect 101 22 103 24
rect 32 10 34 12
rect 80 10 82 12
rect 178 20 180 22
rect 112 10 114 12
rect 226 22 228 24
rect 296 22 298 24
rect 306 22 308 24
rect 196 10 198 12
rect 237 10 239 12
rect 285 10 287 12
rect 383 20 385 22
rect 317 10 319 12
rect 401 10 403 12
rect -194 -2 -192 0
rect -245 -19 -243 -17
rect -110 -2 -108 0
rect -89 -2 -87 0
rect -205 -14 -203 -12
rect -128 -12 -126 -10
rect -5 -2 -3 0
rect -100 -14 -98 -12
rect -23 -12 -21 -10
rect 56 -2 58 0
rect 5 -19 7 -17
rect 140 -2 142 0
rect 161 -2 163 0
rect 45 -14 47 -12
rect 122 -12 124 -10
rect 245 -2 247 0
rect 150 -14 152 -12
rect 227 -12 229 -10
rect 306 -2 308 0
rect 255 -19 257 -17
rect 390 -2 392 0
rect 411 -2 413 0
rect 295 -14 297 -12
rect 372 -12 374 -10
rect 495 -2 497 0
rect 400 -14 402 -12
rect 477 -12 479 -10
rect 556 -2 558 0
rect 505 -19 507 -17
rect 640 -2 642 0
rect 661 -2 663 0
rect 545 -14 547 -12
rect 622 -12 624 -10
rect 745 -2 747 0
rect 650 -14 652 -12
rect 727 -12 729 -10
<< ntiect1 >>
rect 50 82 52 84
rect 90 82 92 84
rect 128 82 130 84
rect 202 82 204 84
rect 255 82 257 84
rect 295 82 297 84
rect 333 82 335 84
rect 407 82 409 84
rect 22 70 24 72
rect 90 70 92 72
rect 102 70 104 72
rect 176 70 178 72
rect 227 70 229 72
rect 295 70 297 72
rect 307 70 309 72
rect 381 70 383 72
rect -244 -62 -242 -60
rect -204 -62 -202 -60
rect -130 -62 -128 -60
rect -99 -62 -97 -60
rect -25 -62 -23 -60
rect 6 -62 8 -60
rect 46 -62 48 -60
rect 120 -62 122 -60
rect 151 -62 153 -60
rect 225 -62 227 -60
rect 256 -62 258 -60
rect 296 -62 298 -60
rect 370 -62 372 -60
rect 401 -62 403 -60
rect 475 -62 477 -60
rect 506 -62 508 -60
rect 546 -62 548 -60
rect 620 -62 622 -60
rect 651 -62 653 -60
rect 725 -62 727 -60
<< ptiect1 >>
rect 50 142 52 144
rect 90 142 92 144
rect 161 142 163 144
rect 202 142 204 144
rect 255 142 257 144
rect 295 142 297 144
rect 366 142 368 144
rect 407 142 409 144
rect 22 10 24 12
rect 90 10 92 12
rect 102 10 104 12
rect 143 10 145 12
rect 227 10 229 12
rect 295 10 297 12
rect 307 10 309 12
rect 348 10 350 12
rect -244 -2 -242 0
rect -204 -2 -202 0
rect -163 -2 -161 0
rect -99 -2 -97 0
rect -58 -2 -56 0
rect 6 -2 8 0
rect 46 -2 48 0
rect 87 -2 89 0
rect 151 -2 153 0
rect 192 -2 194 0
rect 256 -2 258 0
rect 296 -2 298 0
rect 337 -2 339 0
rect 401 -2 403 0
rect 442 -2 444 0
rect 506 -2 508 0
rect 546 -2 548 0
rect 587 -2 589 0
rect 651 -2 653 0
rect 692 -2 694 0
<< pdifct0 >>
rect 21 92 23 94
rect 31 99 33 101
rect 31 92 33 94
rect 41 94 43 96
rect 61 92 63 94
rect 71 99 73 101
rect 71 92 73 94
rect 81 94 83 96
rect 108 91 110 93
rect 128 106 130 108
rect 128 99 130 101
rect 144 92 146 94
rect 144 85 146 87
rect 154 106 156 108
rect 173 92 175 94
rect 183 99 185 101
rect 183 92 185 94
rect 193 94 195 96
rect 226 92 228 94
rect 236 99 238 101
rect 236 92 238 94
rect 246 94 248 96
rect 266 92 268 94
rect 276 99 278 101
rect 276 92 278 94
rect 286 94 288 96
rect 313 91 315 93
rect 333 106 335 108
rect 333 99 335 101
rect 349 92 351 94
rect 349 85 351 87
rect 359 106 361 108
rect 378 92 380 94
rect 388 99 390 101
rect 388 92 390 94
rect 398 94 400 96
rect 31 58 33 60
rect 41 60 43 62
rect 41 53 43 55
rect 51 60 53 62
rect 61 60 63 62
rect 71 60 73 62
rect 71 53 73 55
rect 81 58 83 60
rect 111 58 113 60
rect 121 60 123 62
rect 121 53 123 55
rect 131 60 133 62
rect 150 46 152 48
rect 160 67 162 69
rect 160 60 162 62
rect 176 53 178 55
rect 176 46 178 48
rect 196 61 198 63
rect 236 58 238 60
rect 246 60 248 62
rect 246 53 248 55
rect 256 60 258 62
rect 266 60 268 62
rect 276 60 278 62
rect 276 53 278 55
rect 286 58 288 60
rect 316 58 318 60
rect 326 60 328 62
rect 326 53 328 55
rect 336 60 338 62
rect 355 46 357 48
rect 365 67 367 69
rect 365 60 367 62
rect 381 53 383 55
rect 381 46 383 48
rect 401 61 403 63
rect -234 -59 -232 -57
rect -215 -52 -213 -50
rect -156 -38 -154 -36
rect -195 -50 -193 -48
rect -185 -45 -183 -43
rect -185 -52 -183 -50
rect -175 -52 -173 -50
rect -146 -52 -144 -50
rect -130 -38 -128 -36
rect -130 -45 -128 -43
rect -146 -59 -144 -57
rect -110 -53 -108 -51
rect -51 -38 -49 -36
rect -90 -50 -88 -48
rect -80 -45 -78 -43
rect -80 -52 -78 -50
rect -70 -52 -68 -50
rect -41 -52 -39 -50
rect -25 -38 -23 -36
rect -25 -45 -23 -43
rect -41 -59 -39 -57
rect -5 -53 -3 -51
rect 16 -59 18 -57
rect 35 -52 37 -50
rect 94 -38 96 -36
rect 55 -50 57 -48
rect 65 -45 67 -43
rect 65 -52 67 -50
rect 75 -52 77 -50
rect 104 -52 106 -50
rect 120 -38 122 -36
rect 120 -45 122 -43
rect 104 -59 106 -57
rect 140 -53 142 -51
rect 199 -38 201 -36
rect 160 -50 162 -48
rect 170 -45 172 -43
rect 170 -52 172 -50
rect 180 -52 182 -50
rect 209 -52 211 -50
rect 225 -38 227 -36
rect 225 -45 227 -43
rect 209 -59 211 -57
rect 245 -53 247 -51
rect 266 -59 268 -57
rect 285 -52 287 -50
rect 344 -38 346 -36
rect 305 -50 307 -48
rect 315 -45 317 -43
rect 315 -52 317 -50
rect 325 -52 327 -50
rect 354 -52 356 -50
rect 370 -38 372 -36
rect 370 -45 372 -43
rect 354 -59 356 -57
rect 390 -53 392 -51
rect 449 -38 451 -36
rect 410 -50 412 -48
rect 420 -45 422 -43
rect 420 -52 422 -50
rect 430 -52 432 -50
rect 459 -52 461 -50
rect 475 -38 477 -36
rect 475 -45 477 -43
rect 459 -59 461 -57
rect 495 -53 497 -51
rect 516 -59 518 -57
rect 535 -52 537 -50
rect 594 -38 596 -36
rect 555 -50 557 -48
rect 565 -45 567 -43
rect 565 -52 567 -50
rect 575 -52 577 -50
rect 604 -52 606 -50
rect 620 -38 622 -36
rect 620 -45 622 -43
rect 604 -59 606 -57
rect 640 -53 642 -51
rect 699 -38 701 -36
rect 660 -50 662 -48
rect 670 -45 672 -43
rect 670 -52 672 -50
rect 680 -52 682 -50
rect 709 -52 711 -50
rect 725 -38 727 -36
rect 725 -45 727 -43
rect 709 -59 711 -57
rect 745 -53 747 -51
<< pdifct1 >>
rect 51 106 53 108
rect 51 99 53 101
rect 91 106 93 108
rect 91 99 93 101
rect 118 99 120 101
rect 203 106 205 108
rect 203 99 205 101
rect 256 106 258 108
rect 256 99 258 101
rect 296 106 298 108
rect 296 99 298 101
rect 323 99 325 101
rect 408 106 410 108
rect 408 99 410 101
rect 21 53 23 55
rect 21 46 23 48
rect 91 53 93 55
rect 91 46 93 48
rect 101 53 103 55
rect 101 46 103 48
rect 186 53 188 55
rect 226 53 228 55
rect 226 46 228 48
rect 296 53 298 55
rect 296 46 298 48
rect 306 53 308 55
rect 306 46 308 48
rect 391 53 393 55
rect -245 -42 -243 -40
rect -245 -49 -243 -47
rect -205 -38 -203 -36
rect -205 -45 -203 -43
rect -120 -45 -118 -43
rect -100 -38 -98 -36
rect -100 -45 -98 -43
rect -15 -45 -13 -43
rect 5 -42 7 -40
rect 5 -49 7 -47
rect 45 -38 47 -36
rect 45 -45 47 -43
rect 130 -45 132 -43
rect 150 -38 152 -36
rect 150 -45 152 -43
rect 235 -45 237 -43
rect 255 -42 257 -40
rect 255 -49 257 -47
rect 295 -38 297 -36
rect 295 -45 297 -43
rect 380 -45 382 -43
rect 400 -38 402 -36
rect 400 -45 402 -43
rect 485 -45 487 -43
rect 505 -42 507 -40
rect 505 -49 507 -47
rect 545 -38 547 -36
rect 545 -45 547 -43
rect 630 -45 632 -43
rect 650 -38 652 -36
rect 650 -45 652 -43
rect 735 -45 737 -43
<< alu0 >>
rect 19 134 39 135
rect 19 132 21 134
rect 23 132 39 134
rect 19 131 39 132
rect 35 127 39 131
rect 59 134 79 135
rect 59 132 61 134
rect 63 132 79 134
rect 59 131 79 132
rect 50 128 51 130
rect 35 123 47 127
rect 43 118 47 123
rect 43 116 44 118
rect 46 116 47 118
rect 43 104 47 116
rect 75 127 79 131
rect 146 135 152 141
rect 90 128 91 130
rect 75 123 87 127
rect 83 118 87 123
rect 83 116 84 118
rect 86 116 87 118
rect 30 101 47 104
rect 30 99 31 101
rect 33 100 47 101
rect 33 99 34 100
rect 19 94 25 95
rect 19 92 21 94
rect 23 92 25 94
rect 19 85 25 92
rect 30 94 34 99
rect 83 104 87 116
rect 70 101 87 104
rect 70 99 71 101
rect 73 100 87 101
rect 73 99 74 100
rect 30 92 31 94
rect 33 92 34 94
rect 30 90 34 92
rect 39 96 45 97
rect 39 94 41 96
rect 43 94 45 96
rect 39 85 45 94
rect 59 94 65 95
rect 59 92 61 94
rect 63 92 65 94
rect 59 85 65 92
rect 70 94 74 99
rect 135 132 139 134
rect 146 133 148 135
rect 150 133 152 135
rect 146 132 152 133
rect 171 134 191 135
rect 171 132 173 134
rect 175 132 191 134
rect 135 130 136 132
rect 138 130 139 132
rect 171 131 191 132
rect 135 127 139 130
rect 115 123 139 127
rect 115 119 119 123
rect 161 127 165 129
rect 161 125 162 127
rect 164 125 165 127
rect 114 117 119 119
rect 114 115 115 117
rect 117 115 119 117
rect 123 118 139 119
rect 123 116 125 118
rect 127 116 139 118
rect 123 115 139 116
rect 114 113 119 115
rect 115 111 119 113
rect 115 108 131 111
rect 115 107 128 108
rect 127 106 128 107
rect 130 106 131 108
rect 127 101 131 106
rect 127 99 128 101
rect 130 99 131 101
rect 127 97 131 99
rect 135 109 139 115
rect 161 119 165 125
rect 154 115 165 119
rect 187 127 191 131
rect 224 134 244 135
rect 224 132 226 134
rect 228 132 244 134
rect 224 131 244 132
rect 202 128 203 130
rect 187 123 199 127
rect 195 118 199 123
rect 195 116 196 118
rect 198 116 199 118
rect 154 109 158 115
rect 135 108 158 109
rect 135 106 154 108
rect 156 106 158 108
rect 135 105 158 106
rect 70 92 71 94
rect 73 92 74 94
rect 70 90 74 92
rect 79 96 85 97
rect 79 94 81 96
rect 83 94 85 96
rect 135 94 139 105
rect 195 104 199 116
rect 240 127 244 131
rect 264 134 284 135
rect 264 132 266 134
rect 268 132 284 134
rect 264 131 284 132
rect 255 128 256 130
rect 240 123 252 127
rect 248 118 252 123
rect 248 116 249 118
rect 251 116 252 118
rect 182 101 199 104
rect 182 99 183 101
rect 185 100 199 101
rect 185 99 186 100
rect 79 85 85 94
rect 106 93 139 94
rect 106 91 108 93
rect 110 91 139 93
rect 106 90 139 91
rect 143 94 147 96
rect 143 92 144 94
rect 146 92 147 94
rect 143 87 147 92
rect 171 94 177 95
rect 171 92 173 94
rect 175 92 177 94
rect 143 85 144 87
rect 146 85 147 87
rect 171 85 177 92
rect 182 94 186 99
rect 248 104 252 116
rect 280 127 284 131
rect 351 135 357 141
rect 295 128 296 130
rect 280 123 292 127
rect 288 118 292 123
rect 288 116 289 118
rect 291 116 292 118
rect 235 101 252 104
rect 235 99 236 101
rect 238 100 252 101
rect 238 99 239 100
rect 182 92 183 94
rect 185 92 186 94
rect 182 90 186 92
rect 191 96 197 97
rect 191 94 193 96
rect 195 94 197 96
rect 191 85 197 94
rect 224 94 230 95
rect 224 92 226 94
rect 228 92 230 94
rect 224 85 230 92
rect 235 94 239 99
rect 288 104 292 116
rect 275 101 292 104
rect 275 99 276 101
rect 278 100 292 101
rect 278 99 279 100
rect 235 92 236 94
rect 238 92 239 94
rect 235 90 239 92
rect 244 96 250 97
rect 244 94 246 96
rect 248 94 250 96
rect 244 85 250 94
rect 264 94 270 95
rect 264 92 266 94
rect 268 92 270 94
rect 264 85 270 92
rect 275 94 279 99
rect 340 132 344 134
rect 351 133 353 135
rect 355 133 357 135
rect 351 132 357 133
rect 376 134 396 135
rect 376 132 378 134
rect 380 132 396 134
rect 340 130 341 132
rect 343 130 344 132
rect 376 131 396 132
rect 340 127 344 130
rect 320 123 344 127
rect 320 119 324 123
rect 366 127 370 129
rect 366 125 367 127
rect 369 125 370 127
rect 319 117 324 119
rect 319 115 320 117
rect 322 115 324 117
rect 328 118 344 119
rect 328 116 330 118
rect 332 116 344 118
rect 328 115 344 116
rect 319 113 324 115
rect 320 111 324 113
rect 320 108 336 111
rect 320 107 333 108
rect 332 106 333 107
rect 335 106 336 108
rect 332 101 336 106
rect 332 99 333 101
rect 335 99 336 101
rect 332 97 336 99
rect 340 109 344 115
rect 366 119 370 125
rect 359 115 370 119
rect 392 127 396 131
rect 407 128 408 130
rect 392 123 404 127
rect 400 118 404 123
rect 400 116 401 118
rect 403 116 404 118
rect 359 109 363 115
rect 340 108 363 109
rect 340 106 359 108
rect 361 106 363 108
rect 340 105 363 106
rect 275 92 276 94
rect 278 92 279 94
rect 275 90 279 92
rect 284 96 290 97
rect 284 94 286 96
rect 288 94 290 96
rect 340 94 344 105
rect 400 104 404 116
rect 387 101 404 104
rect 387 99 388 101
rect 390 100 404 101
rect 390 99 391 100
rect 284 85 290 94
rect 311 93 344 94
rect 311 91 313 93
rect 315 91 344 93
rect 311 90 344 91
rect 348 94 352 96
rect 348 92 349 94
rect 351 92 352 94
rect 348 87 352 92
rect 376 94 382 95
rect 376 92 378 94
rect 380 92 382 94
rect 348 85 349 87
rect 351 85 352 87
rect 376 85 382 92
rect 387 94 391 99
rect 387 92 388 94
rect 390 92 391 94
rect 387 90 391 92
rect 396 96 402 97
rect 396 94 398 96
rect 400 94 402 96
rect 396 85 402 94
rect 29 60 35 69
rect 29 58 31 60
rect 33 58 35 60
rect 29 57 35 58
rect 40 62 44 64
rect 40 60 41 62
rect 43 60 44 62
rect 40 55 44 60
rect 49 62 55 69
rect 49 60 51 62
rect 53 60 55 62
rect 49 59 55 60
rect 59 62 65 69
rect 59 60 61 62
rect 63 60 65 62
rect 59 59 65 60
rect 70 62 74 64
rect 70 60 71 62
rect 73 60 74 62
rect 40 54 41 55
rect 27 53 41 54
rect 43 53 44 55
rect 27 50 44 53
rect 27 38 31 50
rect 70 55 74 60
rect 79 60 85 69
rect 79 58 81 60
rect 83 58 85 60
rect 79 57 85 58
rect 109 60 115 69
rect 109 58 111 60
rect 113 58 115 60
rect 109 57 115 58
rect 120 62 124 64
rect 120 60 121 62
rect 123 60 124 62
rect 70 53 71 55
rect 73 54 74 55
rect 73 53 87 54
rect 70 50 87 53
rect 27 36 28 38
rect 30 36 31 38
rect 27 31 31 36
rect 27 27 39 31
rect 23 24 24 26
rect 35 23 39 27
rect 83 38 87 50
rect 83 36 84 38
rect 86 36 87 38
rect 83 31 87 36
rect 75 27 87 31
rect 75 23 79 27
rect 90 24 91 26
rect 35 22 55 23
rect 35 20 51 22
rect 53 20 55 22
rect 35 19 55 20
rect 59 22 79 23
rect 59 20 61 22
rect 63 20 79 22
rect 59 19 79 20
rect 120 55 124 60
rect 129 62 135 69
rect 159 67 160 69
rect 162 67 163 69
rect 129 60 131 62
rect 133 60 135 62
rect 129 59 135 60
rect 159 62 163 67
rect 159 60 160 62
rect 162 60 163 62
rect 159 58 163 60
rect 167 63 200 64
rect 167 61 196 63
rect 198 61 200 63
rect 167 60 200 61
rect 234 60 240 69
rect 120 54 121 55
rect 107 53 121 54
rect 123 53 124 55
rect 107 50 124 53
rect 107 38 111 50
rect 167 49 171 60
rect 234 58 236 60
rect 238 58 240 60
rect 234 57 240 58
rect 245 62 249 64
rect 245 60 246 62
rect 248 60 249 62
rect 148 48 171 49
rect 148 46 150 48
rect 152 46 171 48
rect 148 45 171 46
rect 148 39 152 45
rect 107 36 108 38
rect 110 36 111 38
rect 107 31 111 36
rect 107 27 119 31
rect 103 24 104 26
rect 115 23 119 27
rect 141 35 152 39
rect 141 29 145 35
rect 167 39 171 45
rect 175 55 179 57
rect 175 53 176 55
rect 178 53 179 55
rect 175 48 179 53
rect 175 46 176 48
rect 178 47 179 48
rect 178 46 191 47
rect 175 43 191 46
rect 187 41 191 43
rect 187 39 192 41
rect 167 38 183 39
rect 167 36 179 38
rect 181 36 183 38
rect 167 35 183 36
rect 187 37 189 39
rect 191 37 192 39
rect 187 35 192 37
rect 141 27 142 29
rect 144 27 145 29
rect 141 25 145 27
rect 187 31 191 35
rect 167 27 191 31
rect 167 24 171 27
rect 115 22 135 23
rect 167 22 168 24
rect 170 22 171 24
rect 115 20 131 22
rect 133 20 135 22
rect 115 19 135 20
rect 154 21 160 22
rect 154 19 156 21
rect 158 19 160 21
rect 167 20 171 22
rect 245 55 249 60
rect 254 62 260 69
rect 254 60 256 62
rect 258 60 260 62
rect 254 59 260 60
rect 264 62 270 69
rect 264 60 266 62
rect 268 60 270 62
rect 264 59 270 60
rect 275 62 279 64
rect 275 60 276 62
rect 278 60 279 62
rect 245 54 246 55
rect 232 53 246 54
rect 248 53 249 55
rect 232 50 249 53
rect 232 38 236 50
rect 275 55 279 60
rect 284 60 290 69
rect 284 58 286 60
rect 288 58 290 60
rect 284 57 290 58
rect 314 60 320 69
rect 314 58 316 60
rect 318 58 320 60
rect 314 57 320 58
rect 325 62 329 64
rect 325 60 326 62
rect 328 60 329 62
rect 275 53 276 55
rect 278 54 279 55
rect 278 53 292 54
rect 275 50 292 53
rect 232 36 233 38
rect 235 36 236 38
rect 232 31 236 36
rect 232 27 244 31
rect 228 24 229 26
rect 154 13 160 19
rect 240 23 244 27
rect 288 38 292 50
rect 288 36 289 38
rect 291 36 292 38
rect 288 31 292 36
rect 280 27 292 31
rect 280 23 284 27
rect 295 24 296 26
rect 240 22 260 23
rect 240 20 256 22
rect 258 20 260 22
rect 240 19 260 20
rect 264 22 284 23
rect 264 20 266 22
rect 268 20 284 22
rect 264 19 284 20
rect 325 55 329 60
rect 334 62 340 69
rect 364 67 365 69
rect 367 67 368 69
rect 334 60 336 62
rect 338 60 340 62
rect 334 59 340 60
rect 364 62 368 67
rect 364 60 365 62
rect 367 60 368 62
rect 364 58 368 60
rect 372 63 405 64
rect 372 61 401 63
rect 403 61 405 63
rect 372 60 405 61
rect 325 54 326 55
rect 312 53 326 54
rect 328 53 329 55
rect 312 50 329 53
rect 312 38 316 50
rect 372 49 376 60
rect 353 48 376 49
rect 353 46 355 48
rect 357 46 376 48
rect 353 45 376 46
rect 353 39 357 45
rect 312 36 313 38
rect 315 36 316 38
rect 312 31 316 36
rect 312 27 324 31
rect 308 24 309 26
rect 320 23 324 27
rect 346 35 357 39
rect 346 29 350 35
rect 372 39 376 45
rect 380 55 384 57
rect 380 53 381 55
rect 383 53 384 55
rect 380 48 384 53
rect 380 46 381 48
rect 383 47 384 48
rect 383 46 396 47
rect 380 43 396 46
rect 392 41 396 43
rect 392 39 397 41
rect 372 38 388 39
rect 372 36 384 38
rect 386 36 388 38
rect 372 35 388 36
rect 392 37 394 39
rect 396 37 397 39
rect 392 35 397 37
rect 346 27 347 29
rect 349 27 350 29
rect 346 25 350 27
rect 392 31 396 35
rect 372 27 396 31
rect 372 24 376 27
rect 320 22 340 23
rect 372 22 373 24
rect 375 22 376 24
rect 320 20 336 22
rect 338 20 340 22
rect 320 19 340 20
rect 359 21 365 22
rect 359 19 361 21
rect 363 19 365 21
rect 372 20 376 22
rect 359 13 365 19
rect -236 -4 -230 -3
rect -236 -6 -234 -4
rect -232 -6 -230 -4
rect -236 -7 -230 -6
rect -217 -4 -211 -3
rect -217 -6 -215 -4
rect -213 -6 -211 -4
rect -217 -7 -211 -6
rect -152 -9 -146 -3
rect -191 -10 -171 -9
rect -191 -12 -175 -10
rect -173 -12 -171 -10
rect -152 -11 -150 -9
rect -148 -11 -146 -9
rect -152 -12 -146 -11
rect -139 -12 -135 -10
rect -191 -13 -171 -12
rect -239 -17 -221 -16
rect -239 -19 -225 -17
rect -223 -19 -221 -17
rect -239 -20 -221 -19
rect -239 -26 -235 -20
rect -203 -16 -202 -14
rect -191 -17 -187 -13
rect -139 -14 -138 -12
rect -136 -14 -135 -12
rect -239 -28 -238 -26
rect -236 -28 -235 -26
rect -243 -49 -242 -38
rect -239 -41 -235 -28
rect -220 -33 -214 -32
rect -239 -45 -224 -41
rect -228 -49 -224 -45
rect -199 -21 -187 -17
rect -199 -26 -195 -21
rect -199 -28 -198 -26
rect -196 -28 -195 -26
rect -199 -40 -195 -28
rect -165 -17 -161 -15
rect -165 -19 -164 -17
rect -162 -19 -161 -17
rect -165 -25 -161 -19
rect -139 -17 -135 -14
rect -139 -21 -115 -17
rect -165 -29 -154 -25
rect -158 -35 -154 -29
rect -119 -25 -115 -21
rect -139 -26 -123 -25
rect -139 -28 -127 -26
rect -125 -28 -123 -26
rect -139 -29 -123 -28
rect -119 -27 -114 -25
rect -119 -29 -117 -27
rect -115 -29 -114 -27
rect -139 -35 -135 -29
rect -119 -31 -114 -29
rect -119 -33 -115 -31
rect -158 -36 -135 -35
rect -158 -38 -156 -36
rect -154 -38 -135 -36
rect -158 -39 -135 -38
rect -199 -43 -182 -40
rect -199 -44 -185 -43
rect -186 -45 -185 -44
rect -183 -45 -182 -43
rect -197 -48 -191 -47
rect -228 -50 -211 -49
rect -228 -52 -215 -50
rect -213 -52 -211 -50
rect -228 -53 -211 -52
rect -197 -50 -195 -48
rect -193 -50 -191 -48
rect -236 -57 -230 -56
rect -236 -59 -234 -57
rect -232 -59 -230 -57
rect -197 -59 -191 -50
rect -186 -50 -182 -45
rect -186 -52 -185 -50
rect -183 -52 -182 -50
rect -186 -54 -182 -52
rect -177 -50 -171 -49
rect -177 -52 -175 -50
rect -173 -52 -171 -50
rect -177 -59 -171 -52
rect -147 -50 -143 -48
rect -147 -52 -146 -50
rect -144 -52 -143 -50
rect -147 -57 -143 -52
rect -139 -50 -135 -39
rect -131 -36 -115 -33
rect -131 -38 -130 -36
rect -128 -37 -115 -36
rect -128 -38 -127 -37
rect -131 -43 -127 -38
rect -131 -45 -130 -43
rect -128 -45 -127 -43
rect -131 -47 -127 -45
rect -47 -9 -41 -3
rect 14 -4 20 -3
rect 14 -6 16 -4
rect 18 -6 20 -4
rect 14 -7 20 -6
rect 33 -4 39 -3
rect 33 -6 35 -4
rect 37 -6 39 -4
rect 33 -7 39 -6
rect -86 -10 -66 -9
rect -86 -12 -70 -10
rect -68 -12 -66 -10
rect -47 -11 -45 -9
rect -43 -11 -41 -9
rect -47 -12 -41 -11
rect -34 -12 -30 -10
rect -86 -13 -66 -12
rect -98 -16 -97 -14
rect -86 -17 -82 -13
rect -34 -14 -33 -12
rect -31 -14 -30 -12
rect -94 -21 -82 -17
rect -94 -26 -90 -21
rect -94 -28 -93 -26
rect -91 -28 -90 -26
rect -94 -40 -90 -28
rect -60 -17 -56 -15
rect -60 -19 -59 -17
rect -57 -19 -56 -17
rect -60 -25 -56 -19
rect -34 -17 -30 -14
rect -34 -21 -10 -17
rect -60 -29 -49 -25
rect -53 -35 -49 -29
rect -14 -25 -10 -21
rect -34 -26 -18 -25
rect -34 -28 -22 -26
rect -20 -28 -18 -26
rect -34 -29 -18 -28
rect -14 -27 -9 -25
rect -14 -29 -12 -27
rect -10 -29 -9 -27
rect -34 -35 -30 -29
rect -14 -31 -9 -29
rect -14 -33 -10 -31
rect -53 -36 -30 -35
rect -53 -38 -51 -36
rect -49 -38 -30 -36
rect -53 -39 -30 -38
rect -94 -43 -77 -40
rect -94 -44 -80 -43
rect -81 -45 -80 -44
rect -78 -45 -77 -43
rect -92 -48 -86 -47
rect -92 -50 -90 -48
rect -88 -50 -86 -48
rect -139 -51 -106 -50
rect -139 -53 -110 -51
rect -108 -53 -106 -51
rect -139 -54 -106 -53
rect -147 -59 -146 -57
rect -144 -59 -143 -57
rect -92 -59 -86 -50
rect -81 -50 -77 -45
rect -81 -52 -80 -50
rect -78 -52 -77 -50
rect -81 -54 -77 -52
rect -72 -50 -66 -49
rect -72 -52 -70 -50
rect -68 -52 -66 -50
rect -72 -59 -66 -52
rect -42 -50 -38 -48
rect -42 -52 -41 -50
rect -39 -52 -38 -50
rect -42 -57 -38 -52
rect -34 -50 -30 -39
rect -26 -36 -10 -33
rect -26 -38 -25 -36
rect -23 -37 -10 -36
rect -23 -38 -22 -37
rect -26 -43 -22 -38
rect 98 -9 104 -3
rect 59 -10 79 -9
rect 59 -12 75 -10
rect 77 -12 79 -10
rect 98 -11 100 -9
rect 102 -11 104 -9
rect 98 -12 104 -11
rect 111 -12 115 -10
rect 59 -13 79 -12
rect -26 -45 -25 -43
rect -23 -45 -22 -43
rect -26 -47 -22 -45
rect 11 -17 29 -16
rect 11 -19 25 -17
rect 27 -19 29 -17
rect 11 -20 29 -19
rect 11 -26 15 -20
rect 47 -16 48 -14
rect 59 -17 63 -13
rect 111 -14 112 -12
rect 114 -14 115 -12
rect 11 -28 12 -26
rect 14 -28 15 -26
rect 7 -49 8 -38
rect 11 -41 15 -28
rect 30 -33 36 -32
rect 11 -45 26 -41
rect 22 -49 26 -45
rect 51 -21 63 -17
rect 51 -26 55 -21
rect 51 -28 52 -26
rect 54 -28 55 -26
rect 51 -40 55 -28
rect 85 -17 89 -15
rect 85 -19 86 -17
rect 88 -19 89 -17
rect 85 -25 89 -19
rect 111 -17 115 -14
rect 111 -21 135 -17
rect 85 -29 96 -25
rect 92 -35 96 -29
rect 131 -25 135 -21
rect 111 -26 127 -25
rect 111 -28 123 -26
rect 125 -28 127 -26
rect 111 -29 127 -28
rect 131 -27 136 -25
rect 131 -29 133 -27
rect 135 -29 136 -27
rect 111 -35 115 -29
rect 131 -31 136 -29
rect 131 -33 135 -31
rect 92 -36 115 -35
rect 92 -38 94 -36
rect 96 -38 115 -36
rect 92 -39 115 -38
rect 51 -43 68 -40
rect 51 -44 65 -43
rect 64 -45 65 -44
rect 67 -45 68 -43
rect 53 -48 59 -47
rect -34 -51 -1 -50
rect -34 -53 -5 -51
rect -3 -53 -1 -51
rect -34 -54 -1 -53
rect 22 -50 39 -49
rect 22 -52 35 -50
rect 37 -52 39 -50
rect 22 -53 39 -52
rect 53 -50 55 -48
rect 57 -50 59 -48
rect -42 -59 -41 -57
rect -39 -59 -38 -57
rect 14 -57 20 -56
rect 14 -59 16 -57
rect 18 -59 20 -57
rect 53 -59 59 -50
rect 64 -50 68 -45
rect 64 -52 65 -50
rect 67 -52 68 -50
rect 64 -54 68 -52
rect 73 -50 79 -49
rect 73 -52 75 -50
rect 77 -52 79 -50
rect 73 -59 79 -52
rect 103 -50 107 -48
rect 103 -52 104 -50
rect 106 -52 107 -50
rect 103 -57 107 -52
rect 111 -50 115 -39
rect 119 -36 135 -33
rect 119 -38 120 -36
rect 122 -37 135 -36
rect 122 -38 123 -37
rect 119 -43 123 -38
rect 119 -45 120 -43
rect 122 -45 123 -43
rect 119 -47 123 -45
rect 203 -9 209 -3
rect 264 -4 270 -3
rect 264 -6 266 -4
rect 268 -6 270 -4
rect 264 -7 270 -6
rect 283 -4 289 -3
rect 283 -6 285 -4
rect 287 -6 289 -4
rect 283 -7 289 -6
rect 164 -10 184 -9
rect 164 -12 180 -10
rect 182 -12 184 -10
rect 203 -11 205 -9
rect 207 -11 209 -9
rect 203 -12 209 -11
rect 216 -12 220 -10
rect 164 -13 184 -12
rect 152 -16 153 -14
rect 164 -17 168 -13
rect 216 -14 217 -12
rect 219 -14 220 -12
rect 156 -21 168 -17
rect 156 -26 160 -21
rect 156 -28 157 -26
rect 159 -28 160 -26
rect 156 -40 160 -28
rect 190 -17 194 -15
rect 190 -19 191 -17
rect 193 -19 194 -17
rect 190 -25 194 -19
rect 216 -17 220 -14
rect 216 -21 240 -17
rect 190 -29 201 -25
rect 197 -35 201 -29
rect 236 -25 240 -21
rect 216 -26 232 -25
rect 216 -28 228 -26
rect 230 -28 232 -26
rect 216 -29 232 -28
rect 236 -27 241 -25
rect 236 -29 238 -27
rect 240 -29 241 -27
rect 216 -35 220 -29
rect 236 -31 241 -29
rect 236 -33 240 -31
rect 197 -36 220 -35
rect 197 -38 199 -36
rect 201 -38 220 -36
rect 197 -39 220 -38
rect 156 -43 173 -40
rect 156 -44 170 -43
rect 169 -45 170 -44
rect 172 -45 173 -43
rect 158 -48 164 -47
rect 158 -50 160 -48
rect 162 -50 164 -48
rect 111 -51 144 -50
rect 111 -53 140 -51
rect 142 -53 144 -51
rect 111 -54 144 -53
rect 103 -59 104 -57
rect 106 -59 107 -57
rect 158 -59 164 -50
rect 169 -50 173 -45
rect 169 -52 170 -50
rect 172 -52 173 -50
rect 169 -54 173 -52
rect 178 -50 184 -49
rect 178 -52 180 -50
rect 182 -52 184 -50
rect 178 -59 184 -52
rect 208 -50 212 -48
rect 208 -52 209 -50
rect 211 -52 212 -50
rect 208 -57 212 -52
rect 216 -50 220 -39
rect 224 -36 240 -33
rect 224 -38 225 -36
rect 227 -37 240 -36
rect 227 -38 228 -37
rect 224 -43 228 -38
rect 348 -9 354 -3
rect 309 -10 329 -9
rect 309 -12 325 -10
rect 327 -12 329 -10
rect 348 -11 350 -9
rect 352 -11 354 -9
rect 348 -12 354 -11
rect 361 -12 365 -10
rect 309 -13 329 -12
rect 224 -45 225 -43
rect 227 -45 228 -43
rect 224 -47 228 -45
rect 261 -17 279 -16
rect 261 -19 275 -17
rect 277 -19 279 -17
rect 261 -20 279 -19
rect 261 -26 265 -20
rect 297 -16 298 -14
rect 309 -17 313 -13
rect 361 -14 362 -12
rect 364 -14 365 -12
rect 261 -28 262 -26
rect 264 -28 265 -26
rect 257 -49 258 -38
rect 261 -41 265 -28
rect 280 -33 286 -32
rect 261 -45 276 -41
rect 272 -49 276 -45
rect 301 -21 313 -17
rect 301 -26 305 -21
rect 301 -28 302 -26
rect 304 -28 305 -26
rect 301 -40 305 -28
rect 335 -17 339 -15
rect 335 -19 336 -17
rect 338 -19 339 -17
rect 335 -25 339 -19
rect 361 -17 365 -14
rect 361 -21 385 -17
rect 335 -29 346 -25
rect 342 -35 346 -29
rect 381 -25 385 -21
rect 361 -26 377 -25
rect 361 -28 373 -26
rect 375 -28 377 -26
rect 361 -29 377 -28
rect 381 -27 386 -25
rect 381 -29 383 -27
rect 385 -29 386 -27
rect 361 -35 365 -29
rect 381 -31 386 -29
rect 381 -33 385 -31
rect 342 -36 365 -35
rect 342 -38 344 -36
rect 346 -38 365 -36
rect 342 -39 365 -38
rect 301 -43 318 -40
rect 301 -44 315 -43
rect 314 -45 315 -44
rect 317 -45 318 -43
rect 303 -48 309 -47
rect 216 -51 249 -50
rect 216 -53 245 -51
rect 247 -53 249 -51
rect 216 -54 249 -53
rect 272 -50 289 -49
rect 272 -52 285 -50
rect 287 -52 289 -50
rect 272 -53 289 -52
rect 303 -50 305 -48
rect 307 -50 309 -48
rect 208 -59 209 -57
rect 211 -59 212 -57
rect 264 -57 270 -56
rect 264 -59 266 -57
rect 268 -59 270 -57
rect 303 -59 309 -50
rect 314 -50 318 -45
rect 314 -52 315 -50
rect 317 -52 318 -50
rect 314 -54 318 -52
rect 323 -50 329 -49
rect 323 -52 325 -50
rect 327 -52 329 -50
rect 323 -59 329 -52
rect 353 -50 357 -48
rect 353 -52 354 -50
rect 356 -52 357 -50
rect 353 -57 357 -52
rect 361 -50 365 -39
rect 369 -36 385 -33
rect 369 -38 370 -36
rect 372 -37 385 -36
rect 372 -38 373 -37
rect 369 -43 373 -38
rect 369 -45 370 -43
rect 372 -45 373 -43
rect 369 -47 373 -45
rect 453 -9 459 -3
rect 514 -4 520 -3
rect 514 -6 516 -4
rect 518 -6 520 -4
rect 514 -7 520 -6
rect 533 -4 539 -3
rect 533 -6 535 -4
rect 537 -6 539 -4
rect 533 -7 539 -6
rect 414 -10 434 -9
rect 414 -12 430 -10
rect 432 -12 434 -10
rect 453 -11 455 -9
rect 457 -11 459 -9
rect 453 -12 459 -11
rect 466 -12 470 -10
rect 414 -13 434 -12
rect 402 -16 403 -14
rect 414 -17 418 -13
rect 466 -14 467 -12
rect 469 -14 470 -12
rect 406 -21 418 -17
rect 406 -26 410 -21
rect 406 -28 407 -26
rect 409 -28 410 -26
rect 406 -40 410 -28
rect 440 -17 444 -15
rect 440 -19 441 -17
rect 443 -19 444 -17
rect 440 -25 444 -19
rect 466 -17 470 -14
rect 466 -21 490 -17
rect 440 -29 451 -25
rect 447 -35 451 -29
rect 486 -25 490 -21
rect 466 -26 482 -25
rect 466 -28 478 -26
rect 480 -28 482 -26
rect 466 -29 482 -28
rect 486 -27 491 -25
rect 486 -29 488 -27
rect 490 -29 491 -27
rect 466 -35 470 -29
rect 486 -31 491 -29
rect 486 -33 490 -31
rect 447 -36 470 -35
rect 447 -38 449 -36
rect 451 -38 470 -36
rect 447 -39 470 -38
rect 406 -43 423 -40
rect 406 -44 420 -43
rect 419 -45 420 -44
rect 422 -45 423 -43
rect 408 -48 414 -47
rect 408 -50 410 -48
rect 412 -50 414 -48
rect 361 -51 394 -50
rect 361 -53 390 -51
rect 392 -53 394 -51
rect 361 -54 394 -53
rect 353 -59 354 -57
rect 356 -59 357 -57
rect 408 -59 414 -50
rect 419 -50 423 -45
rect 419 -52 420 -50
rect 422 -52 423 -50
rect 419 -54 423 -52
rect 428 -50 434 -49
rect 428 -52 430 -50
rect 432 -52 434 -50
rect 428 -59 434 -52
rect 458 -50 462 -48
rect 458 -52 459 -50
rect 461 -52 462 -50
rect 458 -57 462 -52
rect 466 -50 470 -39
rect 474 -36 490 -33
rect 474 -38 475 -36
rect 477 -37 490 -36
rect 477 -38 478 -37
rect 474 -43 478 -38
rect 598 -9 604 -3
rect 559 -10 579 -9
rect 559 -12 575 -10
rect 577 -12 579 -10
rect 598 -11 600 -9
rect 602 -11 604 -9
rect 598 -12 604 -11
rect 611 -12 615 -10
rect 559 -13 579 -12
rect 474 -45 475 -43
rect 477 -45 478 -43
rect 474 -47 478 -45
rect 511 -17 529 -16
rect 511 -19 525 -17
rect 527 -19 529 -17
rect 511 -20 529 -19
rect 511 -26 515 -20
rect 547 -16 548 -14
rect 559 -17 563 -13
rect 611 -14 612 -12
rect 614 -14 615 -12
rect 511 -28 512 -26
rect 514 -28 515 -26
rect 507 -49 508 -38
rect 511 -41 515 -28
rect 530 -33 536 -32
rect 511 -45 526 -41
rect 522 -49 526 -45
rect 551 -21 563 -17
rect 551 -26 555 -21
rect 551 -28 552 -26
rect 554 -28 555 -26
rect 551 -40 555 -28
rect 585 -17 589 -15
rect 585 -19 586 -17
rect 588 -19 589 -17
rect 585 -25 589 -19
rect 611 -17 615 -14
rect 611 -21 635 -17
rect 585 -29 596 -25
rect 592 -35 596 -29
rect 631 -25 635 -21
rect 611 -26 627 -25
rect 611 -28 623 -26
rect 625 -28 627 -26
rect 611 -29 627 -28
rect 631 -27 636 -25
rect 631 -29 633 -27
rect 635 -29 636 -27
rect 611 -35 615 -29
rect 631 -31 636 -29
rect 631 -33 635 -31
rect 592 -36 615 -35
rect 592 -38 594 -36
rect 596 -38 615 -36
rect 592 -39 615 -38
rect 551 -43 568 -40
rect 551 -44 565 -43
rect 564 -45 565 -44
rect 567 -45 568 -43
rect 553 -48 559 -47
rect 466 -51 499 -50
rect 466 -53 495 -51
rect 497 -53 499 -51
rect 466 -54 499 -53
rect 522 -50 539 -49
rect 522 -52 535 -50
rect 537 -52 539 -50
rect 522 -53 539 -52
rect 553 -50 555 -48
rect 557 -50 559 -48
rect 458 -59 459 -57
rect 461 -59 462 -57
rect 514 -57 520 -56
rect 514 -59 516 -57
rect 518 -59 520 -57
rect 553 -59 559 -50
rect 564 -50 568 -45
rect 564 -52 565 -50
rect 567 -52 568 -50
rect 564 -54 568 -52
rect 573 -50 579 -49
rect 573 -52 575 -50
rect 577 -52 579 -50
rect 573 -59 579 -52
rect 603 -50 607 -48
rect 603 -52 604 -50
rect 606 -52 607 -50
rect 603 -57 607 -52
rect 611 -50 615 -39
rect 619 -36 635 -33
rect 619 -38 620 -36
rect 622 -37 635 -36
rect 622 -38 623 -37
rect 619 -43 623 -38
rect 619 -45 620 -43
rect 622 -45 623 -43
rect 619 -47 623 -45
rect 703 -9 709 -3
rect 664 -10 684 -9
rect 664 -12 680 -10
rect 682 -12 684 -10
rect 703 -11 705 -9
rect 707 -11 709 -9
rect 703 -12 709 -11
rect 716 -12 720 -10
rect 664 -13 684 -12
rect 652 -16 653 -14
rect 664 -17 668 -13
rect 716 -14 717 -12
rect 719 -14 720 -12
rect 656 -21 668 -17
rect 656 -26 660 -21
rect 656 -28 657 -26
rect 659 -28 660 -26
rect 656 -40 660 -28
rect 690 -17 694 -15
rect 690 -19 691 -17
rect 693 -19 694 -17
rect 690 -25 694 -19
rect 716 -17 720 -14
rect 716 -21 740 -17
rect 690 -29 701 -25
rect 697 -35 701 -29
rect 736 -25 740 -21
rect 716 -26 732 -25
rect 716 -28 728 -26
rect 730 -28 732 -26
rect 716 -29 732 -28
rect 736 -27 741 -25
rect 736 -29 738 -27
rect 740 -29 741 -27
rect 716 -35 720 -29
rect 736 -31 741 -29
rect 736 -33 740 -31
rect 697 -36 720 -35
rect 697 -38 699 -36
rect 701 -38 720 -36
rect 697 -39 720 -38
rect 656 -43 673 -40
rect 656 -44 670 -43
rect 669 -45 670 -44
rect 672 -45 673 -43
rect 658 -48 664 -47
rect 658 -50 660 -48
rect 662 -50 664 -48
rect 611 -51 644 -50
rect 611 -53 640 -51
rect 642 -53 644 -51
rect 611 -54 644 -53
rect 603 -59 604 -57
rect 606 -59 607 -57
rect 658 -59 664 -50
rect 669 -50 673 -45
rect 669 -52 670 -50
rect 672 -52 673 -50
rect 669 -54 673 -52
rect 678 -50 684 -49
rect 678 -52 680 -50
rect 682 -52 684 -50
rect 678 -59 684 -52
rect 708 -50 712 -48
rect 708 -52 709 -50
rect 711 -52 712 -50
rect 708 -57 712 -52
rect 716 -50 720 -39
rect 724 -36 740 -33
rect 724 -38 725 -36
rect 727 -37 740 -36
rect 727 -38 728 -37
rect 724 -43 728 -38
rect 724 -45 725 -43
rect 727 -45 728 -43
rect 724 -47 728 -45
rect 716 -51 749 -50
rect 716 -53 745 -51
rect 747 -53 749 -51
rect 716 -54 749 -53
rect 708 -59 709 -57
rect 711 -59 712 -57
<< via1 >>
rect 37 116 39 118
rect 52 125 54 127
rect 77 116 79 118
rect 20 100 22 102
rect 60 101 62 103
rect 91 102 93 104
rect 153 125 155 127
rect 180 125 182 127
rect 242 116 244 118
rect 204 113 206 115
rect 172 102 174 104
rect 257 125 259 127
rect 282 116 284 118
rect 225 100 227 102
rect 265 101 267 103
rect 296 102 298 104
rect 358 125 360 127
rect 385 125 387 127
rect 409 113 411 115
rect 377 102 379 104
rect 52 53 54 55
rect 60 44 62 46
rect 35 36 37 38
rect 77 36 79 38
rect 92 27 94 29
rect 148 60 150 62
rect 124 27 126 29
rect 151 27 153 29
rect 257 53 259 55
rect 265 44 267 46
rect 240 36 242 38
rect 282 36 284 38
rect 297 27 299 29
rect 353 60 355 62
rect 329 27 331 29
rect 356 27 358 29
rect -214 -45 -212 -43
rect -182 -19 -180 -17
rect -155 -19 -153 -17
rect -109 -19 -107 -17
rect -77 -19 -75 -17
rect -100 -45 -98 -43
rect -50 -19 -48 -17
rect -67 -37 -65 -35
rect 4 -37 6 -35
rect 36 -45 38 -43
rect 68 -19 70 -17
rect 95 -19 97 -17
rect 141 -19 143 -17
rect 173 -19 175 -17
rect 150 -45 152 -43
rect 200 -19 202 -17
rect 185 -37 187 -35
rect 254 -37 256 -35
rect 286 -45 288 -43
rect 318 -19 320 -17
rect 345 -19 347 -17
rect 391 -19 393 -17
rect 423 -19 425 -17
rect 400 -45 402 -43
rect 450 -19 452 -17
rect 435 -37 437 -35
rect 504 -37 506 -35
rect 536 -45 538 -43
rect 568 -19 570 -17
rect 595 -19 597 -17
rect 641 -19 643 -17
rect 673 -19 675 -17
rect 650 -45 652 -43
rect 700 -19 702 -17
<< labels >>
rlabel alu1 141 73 141 73 1 Vdd
rlabel alu1 117 73 117 73 6 vdd
rlabel alu1 139 8 139 8 1 Vss
rlabel alu1 37 9 37 9 6 vss
rlabel alu1 37 73 37 73 6 vdd
rlabel alu1 77 9 77 9 4 vss
rlabel alu1 77 73 77 73 4 vdd
rlabel alu1 167 146 167 146 5 Vss
rlabel alu1 189 81 189 81 2 vdd
rlabel alu1 165 81 165 81 5 Vdd
rlabel alu1 37 81 37 81 2 vdd
rlabel alu1 37 145 37 145 2 vss
rlabel alu1 77 145 77 145 2 vss
rlabel alu1 77 81 77 81 2 vdd
rlabel alu1 234 123 234 123 1 a0
rlabel alu1 274 121 274 121 1 a1
rlabel alu1 282 81 282 81 2 vdd
rlabel alu1 282 145 282 145 2 vss
rlabel alu1 242 145 242 145 2 vss
rlabel alu1 242 81 242 81 2 vdd
rlabel alu1 370 81 370 81 5 Vdd
rlabel alu1 394 81 394 81 2 vdd
rlabel alu1 372 146 372 146 5 Vss
rlabel alu1 282 73 282 73 4 vdd
rlabel alu1 282 9 282 9 4 vss
rlabel alu1 274 32 274 32 1 a1
rlabel alu1 250 31 250 31 1 a0
rlabel alu1 242 73 242 73 6 vdd
rlabel alu1 242 9 242 9 6 vss
rlabel alu1 344 8 344 8 1 Vss
rlabel alu1 322 73 322 73 6 vdd
rlabel alu1 346 73 346 73 1 Vdd
rlabel alu1 306 35 306 35 1 p13
rlabel alu1 226 37 226 37 1 p10
rlabel alu1 403 40 403 40 1 p12
rlabel alu1 313 114 313 114 1 p11
rlabel alu1 21 37 21 37 1 p20
rlabel alu1 101 35 101 35 1 p23
rlabel alu1 198 40 198 40 1 p22
rlabel alu1 -165 -63 -165 -63 5 Vdd
rlabel alu1 -189 -63 -189 -63 8 vdd
rlabel alu1 -167 2 -167 2 5 Vss
rlabel alu1 -60 -63 -60 -63 5 Vdd
rlabel alu1 -84 -63 -84 -63 8 vdd
rlabel alu1 -62 2 -62 2 5 Vss
rlabel alu1 -229 -63 -229 -63 8 vdd
rlabel alu1 85 -63 85 -63 5 Vdd
rlabel alu1 61 -63 61 -63 8 vdd
rlabel alu1 83 2 83 2 5 Vss
rlabel alu1 190 -63 190 -63 5 Vdd
rlabel alu1 166 -63 166 -63 8 vdd
rlabel alu1 188 2 188 2 5 Vss
rlabel alu1 21 -63 21 -63 8 vdd
rlabel alu1 271 -63 271 -63 8 vdd
rlabel alu1 438 2 438 2 5 Vss
rlabel alu1 416 -63 416 -63 8 vdd
rlabel alu1 440 -63 440 -63 5 Vdd
rlabel alu1 333 2 333 2 5 Vss
rlabel alu1 311 -63 311 -63 8 vdd
rlabel alu1 335 -63 335 -63 5 Vdd
rlabel alu1 585 -63 585 -63 5 Vdd
rlabel alu1 561 -63 561 -63 8 vdd
rlabel alu1 583 2 583 2 5 Vss
rlabel alu1 690 -63 690 -63 5 Vdd
rlabel alu1 666 -63 666 -63 8 vdd
rlabel alu1 688 2 688 2 5 Vss
rlabel alu1 521 -63 521 -63 8 vdd
rlabel alu1 -156 -51 -156 -51 5 p23
rlabel alu1 -147 -26 -147 -26 5 p13
rlabel alu1 94 -51 94 -51 5 p22
rlabel alu1 103 -26 103 -26 5 p12
rlabel alu1 344 -51 344 -51 5 p21
rlabel alu1 353 -26 353 -26 5 p11
rlabel alu1 594 -51 594 -51 5 p20
rlabel alu1 603 -26 603 -26 5 p10
rlabel via1 258 53 258 53 1 b2
rlabel alu1 266 53 266 53 1 b3
rlabel alu1 274 109 274 109 1 b2
rlabel via1 226 101 226 101 1 b3
rlabel via1 21 101 21 101 1 b1
rlabel alu1 69 109 69 109 1 b0
rlabel via1 53 53 53 53 1 b0
rlabel alu1 61 53 61 53 1 b1
rlabel alu1 45 31 45 31 1 a2
rlabel alu1 69 32 69 32 1 a3
rlabel alu1 29 123 29 123 1 a2
rlabel alu1 69 121 69 121 1 a3
rlabel alu1 108 114 108 114 1 p21
rlabel alu1 682 -43 682 -43 1 Vss
rlabel alu1 -245 -34 -245 -34 1 c0
rlabel alu1 -3 -30 -3 -30 1 s03
rlabel alu1 247 -30 247 -30 1 s02
rlabel alu1 497 -30 497 -30 1 s01
rlabel alu1 747 -30 747 -30 1 s00
<< end >>
