magic
tech scmos
timestamp 1607834672
<< ab >>
rect 88 159 94 164
rect 202 159 208 164
rect 4 15 44 159
rect 53 127 157 159
rect 53 95 93 127
rect 94 95 157 127
rect 46 79 51 95
rect 53 79 157 95
rect 53 47 93 79
rect 94 47 157 79
rect 53 15 157 47
rect 167 127 271 159
rect 272 151 276 159
rect 167 114 207 127
rect 208 114 271 127
rect 167 105 271 114
rect 167 95 207 105
rect 208 95 271 105
rect 167 79 271 95
rect 272 79 274 95
rect 167 47 207 79
rect 208 47 271 79
rect 167 15 271 47
rect 272 15 276 23
rect 278 15 318 159
rect 319 151 383 159
rect 322 95 383 151
rect 319 79 383 95
rect 322 23 383 79
rect 319 15 383 23
rect 387 15 451 159
rect 455 15 518 159
rect 520 151 560 159
rect 562 151 632 159
rect 521 95 560 151
rect 563 95 626 151
rect 520 79 560 95
rect 561 79 626 95
rect 627 79 632 95
rect 521 23 560 79
rect 563 23 626 79
rect 520 15 560 23
rect 562 15 632 23
rect 88 10 94 15
rect 202 10 208 15
<< nwell >>
rect -1 47 632 127
<< pwell >>
rect -1 127 632 164
rect -1 10 632 47
<< poly >>
rect 13 142 15 147
rect 23 139 25 144
rect 33 139 35 144
rect 62 144 64 148
rect 75 146 77 151
rect 82 146 84 151
rect 105 155 130 157
rect 105 147 107 155
rect 118 147 120 151
rect 128 147 130 155
rect 138 150 140 155
rect 145 150 147 155
rect 102 145 107 147
rect 102 142 104 145
rect 13 130 15 133
rect 23 130 25 133
rect 13 128 19 130
rect 13 126 15 128
rect 17 126 19 128
rect 13 124 19 126
rect 23 128 29 130
rect 23 126 25 128
rect 27 126 29 128
rect 23 124 29 126
rect 13 121 15 124
rect 26 114 28 124
rect 33 123 35 133
rect 62 130 64 135
rect 75 130 77 135
rect 62 128 68 130
rect 62 126 64 128
rect 66 126 68 128
rect 62 124 68 126
rect 72 128 78 130
rect 72 126 74 128
rect 76 126 78 128
rect 72 124 78 126
rect 33 121 39 123
rect 33 119 35 121
rect 37 119 39 121
rect 62 120 64 124
rect 33 117 39 119
rect 33 114 35 117
rect 13 98 15 103
rect 72 113 74 124
rect 82 122 84 135
rect 176 144 178 148
rect 189 146 191 151
rect 196 146 198 151
rect 219 155 244 157
rect 219 147 221 155
rect 232 147 234 151
rect 242 147 244 155
rect 252 150 254 155
rect 259 150 261 155
rect 118 135 120 138
rect 111 133 120 135
rect 128 134 130 138
rect 138 135 140 138
rect 102 125 104 133
rect 111 131 113 133
rect 115 131 120 133
rect 111 129 120 131
rect 136 133 140 135
rect 136 130 138 133
rect 118 125 120 129
rect 132 128 138 130
rect 145 129 147 138
rect 216 145 221 147
rect 216 142 218 145
rect 176 130 178 135
rect 189 130 191 135
rect 132 126 134 128
rect 136 126 138 128
rect 99 123 112 125
rect 118 123 128 125
rect 132 124 138 126
rect 99 122 101 123
rect 82 120 88 122
rect 82 118 84 120
rect 86 118 88 120
rect 82 116 88 118
rect 95 120 101 122
rect 110 120 112 123
rect 126 120 128 123
rect 136 120 138 124
rect 142 127 148 129
rect 142 125 144 127
rect 146 125 148 127
rect 142 123 148 125
rect 146 120 148 123
rect 176 128 182 130
rect 176 126 178 128
rect 180 126 182 128
rect 176 124 182 126
rect 186 128 192 130
rect 186 126 188 128
rect 190 126 192 128
rect 186 124 192 126
rect 176 120 178 124
rect 95 118 97 120
rect 99 118 101 120
rect 95 116 101 118
rect 82 113 84 116
rect 62 98 64 102
rect 72 95 74 100
rect 82 95 84 100
rect 26 89 28 93
rect 33 89 35 93
rect 126 98 128 102
rect 136 98 138 102
rect 110 89 112 93
rect 186 113 188 124
rect 196 122 198 135
rect 287 146 289 151
rect 294 146 296 151
rect 329 155 348 157
rect 232 135 234 138
rect 225 133 234 135
rect 242 134 244 138
rect 252 135 254 138
rect 216 125 218 133
rect 225 131 227 133
rect 229 131 234 133
rect 225 129 234 131
rect 250 133 254 135
rect 250 130 252 133
rect 232 125 234 129
rect 246 128 252 130
rect 259 129 261 138
rect 307 144 309 148
rect 329 145 331 155
rect 339 147 341 151
rect 346 147 348 155
rect 423 155 442 157
rect 356 147 358 152
rect 363 147 365 152
rect 373 147 375 152
rect 396 147 398 152
rect 406 147 408 152
rect 413 147 415 152
rect 423 147 425 155
rect 430 147 432 151
rect 246 126 248 128
rect 250 126 252 128
rect 213 123 226 125
rect 232 123 242 125
rect 246 124 252 126
rect 213 122 215 123
rect 196 120 202 122
rect 196 118 198 120
rect 200 118 202 120
rect 196 116 202 118
rect 209 120 215 122
rect 224 120 226 123
rect 240 120 242 123
rect 250 120 252 124
rect 256 127 262 129
rect 256 125 258 127
rect 260 125 262 127
rect 256 123 262 125
rect 260 120 262 123
rect 287 122 289 135
rect 294 130 296 135
rect 307 130 309 135
rect 293 128 299 130
rect 293 126 295 128
rect 297 126 299 128
rect 293 124 299 126
rect 303 128 309 130
rect 303 126 305 128
rect 307 126 309 128
rect 303 124 309 126
rect 283 120 289 122
rect 209 118 211 120
rect 213 118 215 120
rect 209 116 215 118
rect 196 113 198 116
rect 176 98 178 102
rect 186 95 188 100
rect 196 95 198 100
rect 146 89 148 93
rect 240 98 242 102
rect 250 98 252 102
rect 224 89 226 93
rect 283 118 285 120
rect 287 118 289 120
rect 283 116 289 118
rect 287 113 289 116
rect 297 113 299 124
rect 307 120 309 124
rect 329 121 331 139
rect 339 130 341 139
rect 335 128 341 130
rect 335 126 337 128
rect 339 126 341 128
rect 335 124 341 126
rect 346 126 348 139
rect 356 136 358 139
rect 352 134 358 136
rect 352 132 354 134
rect 356 132 358 134
rect 352 130 358 132
rect 346 124 358 126
rect 363 125 365 139
rect 440 145 442 155
rect 490 155 509 157
rect 463 147 465 152
rect 473 147 475 152
rect 480 147 482 152
rect 490 147 492 155
rect 497 147 499 151
rect 373 135 375 138
rect 396 135 398 138
rect 370 133 376 135
rect 370 131 372 133
rect 374 131 376 133
rect 370 129 376 131
rect 395 133 401 135
rect 395 131 397 133
rect 399 131 401 133
rect 395 129 401 131
rect 329 110 331 113
rect 322 108 331 110
rect 339 109 341 124
rect 345 118 351 120
rect 345 116 347 118
rect 349 116 351 118
rect 345 114 351 116
rect 346 109 348 114
rect 356 109 358 124
rect 362 123 368 125
rect 362 121 364 123
rect 366 121 368 123
rect 362 119 368 121
rect 363 109 365 119
rect 373 111 375 129
rect 396 111 398 129
rect 406 125 408 139
rect 413 136 415 139
rect 413 134 419 136
rect 413 132 415 134
rect 417 132 419 134
rect 413 130 419 132
rect 423 126 425 139
rect 403 123 409 125
rect 403 121 405 123
rect 407 121 409 123
rect 403 119 409 121
rect 413 124 425 126
rect 430 130 432 139
rect 430 128 436 130
rect 430 126 432 128
rect 434 126 436 128
rect 430 124 436 126
rect 322 106 324 108
rect 326 106 328 108
rect 322 104 328 106
rect 287 95 289 100
rect 297 95 299 100
rect 307 98 309 102
rect 260 89 262 93
rect 406 109 408 119
rect 413 109 415 124
rect 420 118 426 120
rect 420 116 422 118
rect 424 116 426 118
rect 420 114 426 116
rect 423 109 425 114
rect 430 109 432 124
rect 440 121 442 139
rect 507 145 509 155
rect 589 155 614 157
rect 529 142 531 147
rect 463 135 465 138
rect 462 133 468 135
rect 462 131 464 133
rect 466 131 468 133
rect 462 129 468 131
rect 440 110 442 113
rect 463 111 465 129
rect 473 125 475 139
rect 480 136 482 139
rect 480 134 486 136
rect 480 132 482 134
rect 484 132 486 134
rect 480 130 486 132
rect 490 126 492 139
rect 470 123 476 125
rect 470 121 472 123
rect 474 121 476 123
rect 470 119 476 121
rect 480 124 492 126
rect 497 130 499 139
rect 497 128 503 130
rect 497 126 499 128
rect 501 126 503 128
rect 497 124 503 126
rect 440 108 449 110
rect 443 106 445 108
rect 447 106 449 108
rect 443 104 449 106
rect 473 109 475 119
rect 480 109 482 124
rect 487 118 493 120
rect 487 116 489 118
rect 491 116 493 118
rect 487 114 493 116
rect 490 109 492 114
rect 497 109 499 124
rect 507 121 509 139
rect 539 139 541 144
rect 549 139 551 144
rect 572 150 574 155
rect 579 150 581 155
rect 589 147 591 155
rect 599 147 601 151
rect 612 147 614 155
rect 612 145 617 147
rect 615 142 617 145
rect 529 130 531 133
rect 539 130 541 133
rect 529 128 535 130
rect 529 126 531 128
rect 533 126 535 128
rect 529 124 535 126
rect 539 128 545 130
rect 539 126 541 128
rect 543 126 545 128
rect 539 124 545 126
rect 529 121 531 124
rect 507 110 509 113
rect 507 108 516 110
rect 510 106 512 108
rect 514 106 516 108
rect 510 104 516 106
rect 542 114 544 124
rect 549 123 551 133
rect 572 129 574 138
rect 579 135 581 138
rect 579 133 583 135
rect 589 134 591 138
rect 599 135 601 138
rect 581 130 583 133
rect 599 133 608 135
rect 599 131 604 133
rect 606 131 608 133
rect 571 127 577 129
rect 571 125 573 127
rect 575 125 577 127
rect 571 123 577 125
rect 581 128 587 130
rect 581 126 583 128
rect 585 126 587 128
rect 581 124 587 126
rect 599 129 608 131
rect 599 125 601 129
rect 615 125 617 133
rect 549 121 555 123
rect 549 119 551 121
rect 553 119 555 121
rect 571 120 573 123
rect 581 120 583 124
rect 591 123 601 125
rect 607 123 620 125
rect 591 120 593 123
rect 607 120 609 123
rect 618 122 620 123
rect 618 120 624 122
rect 549 117 555 119
rect 549 114 551 117
rect 529 98 531 103
rect 339 89 341 93
rect 346 89 348 93
rect 356 89 358 93
rect 363 89 365 93
rect 373 89 375 93
rect 396 89 398 93
rect 406 89 408 93
rect 413 89 415 93
rect 423 89 425 93
rect 430 89 432 93
rect 463 89 465 93
rect 473 89 475 93
rect 480 89 482 93
rect 490 89 492 93
rect 497 89 499 93
rect 581 98 583 102
rect 591 98 593 102
rect 542 89 544 93
rect 549 89 551 93
rect 571 89 573 93
rect 618 118 620 120
rect 622 118 624 120
rect 618 116 624 118
rect 607 89 609 93
rect 26 81 28 85
rect 33 81 35 85
rect 13 71 15 76
rect 110 81 112 85
rect 62 72 64 76
rect 72 74 74 79
rect 82 74 84 79
rect 13 50 15 53
rect 26 50 28 60
rect 33 57 35 60
rect 33 55 39 57
rect 33 53 35 55
rect 37 53 39 55
rect 33 51 39 53
rect 13 48 19 50
rect 13 46 15 48
rect 17 46 19 48
rect 13 44 19 46
rect 23 48 29 50
rect 23 46 25 48
rect 27 46 29 48
rect 23 44 29 46
rect 13 41 15 44
rect 23 41 25 44
rect 33 41 35 51
rect 62 50 64 54
rect 72 50 74 61
rect 82 58 84 61
rect 82 56 88 58
rect 82 54 84 56
rect 86 54 88 56
rect 82 52 88 54
rect 95 56 101 58
rect 95 54 97 56
rect 99 54 101 56
rect 146 81 148 85
rect 126 72 128 76
rect 136 72 138 76
rect 224 81 226 85
rect 176 72 178 76
rect 186 74 188 79
rect 196 74 198 79
rect 95 52 101 54
rect 62 48 68 50
rect 62 46 64 48
rect 66 46 68 48
rect 62 44 68 46
rect 72 48 78 50
rect 72 46 74 48
rect 76 46 78 48
rect 72 44 78 46
rect 62 39 64 44
rect 75 39 77 44
rect 82 39 84 52
rect 99 51 101 52
rect 110 51 112 54
rect 126 51 128 54
rect 99 49 112 51
rect 118 49 128 51
rect 136 50 138 54
rect 146 51 148 54
rect 102 41 104 49
rect 118 45 120 49
rect 111 43 120 45
rect 132 48 138 50
rect 132 46 134 48
rect 136 46 138 48
rect 132 44 138 46
rect 142 49 148 51
rect 142 47 144 49
rect 146 47 148 49
rect 142 45 148 47
rect 176 50 178 54
rect 186 50 188 61
rect 196 58 198 61
rect 196 56 202 58
rect 196 54 198 56
rect 200 54 202 56
rect 196 52 202 54
rect 209 56 215 58
rect 209 54 211 56
rect 213 54 215 56
rect 260 81 262 85
rect 240 72 242 76
rect 250 72 252 76
rect 339 81 341 85
rect 346 81 348 85
rect 356 81 358 85
rect 363 81 365 85
rect 373 81 375 85
rect 396 81 398 85
rect 406 81 408 85
rect 413 81 415 85
rect 423 81 425 85
rect 430 81 432 85
rect 463 81 465 85
rect 473 81 475 85
rect 480 81 482 85
rect 490 81 492 85
rect 497 81 499 85
rect 287 74 289 79
rect 297 74 299 79
rect 307 72 309 76
rect 287 58 289 61
rect 283 56 289 58
rect 283 54 285 56
rect 287 54 289 56
rect 209 52 215 54
rect 176 48 182 50
rect 176 46 178 48
rect 180 46 182 48
rect 111 41 113 43
rect 115 41 120 43
rect 13 27 15 32
rect 23 30 25 35
rect 33 30 35 35
rect 62 26 64 30
rect 111 39 120 41
rect 136 41 138 44
rect 118 36 120 39
rect 128 36 130 40
rect 136 39 140 41
rect 138 36 140 39
rect 145 36 147 45
rect 176 44 182 46
rect 186 48 192 50
rect 186 46 188 48
rect 190 46 192 48
rect 186 44 192 46
rect 176 39 178 44
rect 189 39 191 44
rect 196 39 198 52
rect 213 51 215 52
rect 224 51 226 54
rect 240 51 242 54
rect 213 49 226 51
rect 232 49 242 51
rect 250 50 252 54
rect 260 51 262 54
rect 283 52 289 54
rect 216 41 218 49
rect 232 45 234 49
rect 225 43 234 45
rect 246 48 252 50
rect 246 46 248 48
rect 250 46 252 48
rect 246 44 252 46
rect 256 49 262 51
rect 256 47 258 49
rect 260 47 262 49
rect 256 45 262 47
rect 225 41 227 43
rect 229 41 234 43
rect 102 29 104 32
rect 75 23 77 28
rect 82 23 84 28
rect 102 27 107 29
rect 105 19 107 27
rect 118 23 120 27
rect 128 19 130 27
rect 176 26 178 30
rect 225 39 234 41
rect 250 41 252 44
rect 232 36 234 39
rect 242 36 244 40
rect 250 39 254 41
rect 252 36 254 39
rect 259 36 261 45
rect 287 39 289 52
rect 297 50 299 61
rect 322 68 328 70
rect 322 66 324 68
rect 326 66 328 68
rect 322 64 331 66
rect 329 61 331 64
rect 307 50 309 54
rect 293 48 299 50
rect 293 46 295 48
rect 297 46 299 48
rect 293 44 299 46
rect 303 48 309 50
rect 303 46 305 48
rect 307 46 309 48
rect 303 44 309 46
rect 294 39 296 44
rect 307 39 309 44
rect 216 29 218 32
rect 138 19 140 24
rect 145 19 147 24
rect 105 17 130 19
rect 189 23 191 28
rect 196 23 198 28
rect 216 27 221 29
rect 219 19 221 27
rect 232 23 234 27
rect 242 19 244 27
rect 329 35 331 53
rect 339 50 341 65
rect 346 60 348 65
rect 345 58 351 60
rect 345 56 347 58
rect 349 56 351 58
rect 345 54 351 56
rect 356 50 358 65
rect 363 55 365 65
rect 443 68 449 70
rect 443 66 445 68
rect 447 66 449 68
rect 335 48 341 50
rect 335 46 337 48
rect 339 46 341 48
rect 335 44 341 46
rect 339 35 341 44
rect 346 48 358 50
rect 362 53 368 55
rect 362 51 364 53
rect 366 51 368 53
rect 362 49 368 51
rect 346 35 348 48
rect 352 42 358 44
rect 352 40 354 42
rect 356 40 358 42
rect 352 38 358 40
rect 356 35 358 38
rect 363 35 365 49
rect 373 45 375 63
rect 396 45 398 63
rect 406 55 408 65
rect 403 53 409 55
rect 403 51 405 53
rect 407 51 409 53
rect 403 49 409 51
rect 413 50 415 65
rect 423 60 425 65
rect 420 58 426 60
rect 420 56 422 58
rect 424 56 426 58
rect 420 54 426 56
rect 430 50 432 65
rect 440 64 449 66
rect 440 61 442 64
rect 542 81 544 85
rect 549 81 551 85
rect 571 81 573 85
rect 529 71 531 76
rect 510 68 516 70
rect 510 66 512 68
rect 514 66 516 68
rect 370 43 376 45
rect 370 41 372 43
rect 374 41 376 43
rect 370 39 376 41
rect 395 43 401 45
rect 395 41 397 43
rect 399 41 401 43
rect 395 39 401 41
rect 373 36 375 39
rect 396 36 398 39
rect 252 19 254 24
rect 259 19 261 24
rect 287 23 289 28
rect 294 23 296 28
rect 219 17 244 19
rect 307 26 309 30
rect 329 19 331 29
rect 406 35 408 49
rect 413 48 425 50
rect 413 42 419 44
rect 413 40 415 42
rect 417 40 419 42
rect 413 38 419 40
rect 413 35 415 38
rect 423 35 425 48
rect 430 48 436 50
rect 430 46 432 48
rect 434 46 436 48
rect 430 44 436 46
rect 430 35 432 44
rect 440 35 442 53
rect 463 45 465 63
rect 473 55 475 65
rect 470 53 476 55
rect 470 51 472 53
rect 474 51 476 53
rect 470 49 476 51
rect 480 50 482 65
rect 490 60 492 65
rect 487 58 493 60
rect 487 56 489 58
rect 491 56 493 58
rect 487 54 493 56
rect 497 50 499 65
rect 507 64 516 66
rect 507 61 509 64
rect 462 43 468 45
rect 462 41 464 43
rect 466 41 468 43
rect 462 39 468 41
rect 463 36 465 39
rect 339 23 341 27
rect 346 19 348 27
rect 356 22 358 27
rect 363 22 365 27
rect 373 22 375 27
rect 396 22 398 27
rect 406 22 408 27
rect 413 22 415 27
rect 329 17 348 19
rect 423 19 425 27
rect 430 23 432 27
rect 440 19 442 29
rect 473 35 475 49
rect 480 48 492 50
rect 480 42 486 44
rect 480 40 482 42
rect 484 40 486 42
rect 480 38 486 40
rect 480 35 482 38
rect 490 35 492 48
rect 497 48 503 50
rect 497 46 499 48
rect 501 46 503 48
rect 497 44 503 46
rect 497 35 499 44
rect 507 35 509 53
rect 529 50 531 53
rect 542 50 544 60
rect 549 57 551 60
rect 549 55 555 57
rect 549 53 551 55
rect 553 53 555 55
rect 607 81 609 85
rect 581 72 583 76
rect 591 72 593 76
rect 618 56 624 58
rect 618 54 620 56
rect 622 54 624 56
rect 549 51 555 53
rect 571 51 573 54
rect 529 48 535 50
rect 529 46 531 48
rect 533 46 535 48
rect 529 44 535 46
rect 539 48 545 50
rect 539 46 541 48
rect 543 46 545 48
rect 539 44 545 46
rect 529 41 531 44
rect 539 41 541 44
rect 549 41 551 51
rect 571 49 577 51
rect 571 47 573 49
rect 575 47 577 49
rect 571 45 577 47
rect 581 50 583 54
rect 591 51 593 54
rect 607 51 609 54
rect 618 52 624 54
rect 618 51 620 52
rect 581 48 587 50
rect 591 49 601 51
rect 607 49 620 51
rect 581 46 583 48
rect 585 46 587 48
rect 572 36 574 45
rect 581 44 587 46
rect 599 45 601 49
rect 581 41 583 44
rect 579 39 583 41
rect 599 43 608 45
rect 599 41 604 43
rect 606 41 608 43
rect 615 41 617 49
rect 579 36 581 39
rect 589 36 591 40
rect 599 39 608 41
rect 599 36 601 39
rect 463 22 465 27
rect 473 22 475 27
rect 480 22 482 27
rect 423 17 442 19
rect 490 19 492 27
rect 497 23 499 27
rect 507 19 509 29
rect 529 27 531 32
rect 539 30 541 35
rect 549 30 551 35
rect 490 17 509 19
rect 615 29 617 32
rect 612 27 617 29
rect 572 19 574 24
rect 579 19 581 24
rect 589 19 591 27
rect 599 23 601 27
rect 612 19 614 27
rect 589 17 614 19
<< ndif >>
rect 17 150 23 152
rect 17 148 19 150
rect 21 148 23 150
rect 17 146 23 148
rect 36 150 42 152
rect 66 154 73 156
rect 66 152 68 154
rect 70 152 73 154
rect 36 148 38 150
rect 40 148 42 150
rect 36 146 42 148
rect 17 142 21 146
rect 8 139 13 142
rect 6 137 13 139
rect 6 135 8 137
rect 10 135 13 137
rect 6 133 13 135
rect 15 139 21 142
rect 37 139 42 146
rect 66 146 73 152
rect 149 154 155 156
rect 149 152 151 154
rect 153 152 155 154
rect 149 150 155 152
rect 180 154 187 156
rect 180 152 182 154
rect 184 152 187 154
rect 133 147 138 150
rect 66 144 75 146
rect 15 133 23 139
rect 25 137 33 139
rect 25 135 28 137
rect 30 135 33 137
rect 25 133 33 135
rect 35 133 42 139
rect 55 142 62 144
rect 55 140 57 142
rect 59 140 62 142
rect 55 138 62 140
rect 57 135 62 138
rect 64 135 75 144
rect 77 135 82 146
rect 84 144 91 146
rect 84 142 87 144
rect 89 142 91 144
rect 109 145 118 147
rect 109 143 111 145
rect 113 143 118 145
rect 109 142 118 143
rect 84 140 91 142
rect 84 135 89 140
rect 97 139 102 142
rect 95 137 102 139
rect 95 135 97 137
rect 99 135 102 137
rect 95 133 102 135
rect 104 138 118 142
rect 120 142 128 147
rect 120 140 123 142
rect 125 140 128 142
rect 120 138 128 140
rect 130 144 138 147
rect 130 142 133 144
rect 135 142 138 144
rect 130 138 138 142
rect 140 138 145 150
rect 147 138 155 150
rect 180 146 187 152
rect 263 154 269 156
rect 263 152 265 154
rect 267 152 269 154
rect 263 150 269 152
rect 298 154 305 156
rect 298 152 301 154
rect 303 152 305 154
rect 247 147 252 150
rect 180 144 189 146
rect 169 142 176 144
rect 169 140 171 142
rect 173 140 176 142
rect 169 138 176 140
rect 104 133 109 138
rect 171 135 176 138
rect 178 135 189 144
rect 191 135 196 146
rect 198 144 205 146
rect 198 142 201 144
rect 203 142 205 144
rect 223 145 232 147
rect 223 143 225 145
rect 227 143 232 145
rect 223 142 232 143
rect 198 140 205 142
rect 198 135 203 140
rect 211 139 216 142
rect 209 137 216 139
rect 209 135 211 137
rect 213 135 216 137
rect 209 133 216 135
rect 218 138 232 142
rect 234 142 242 147
rect 234 140 237 142
rect 239 140 242 142
rect 234 138 242 140
rect 244 144 252 147
rect 244 142 247 144
rect 249 142 252 144
rect 244 138 252 142
rect 254 138 259 150
rect 261 138 269 150
rect 298 146 305 152
rect 280 144 287 146
rect 280 142 282 144
rect 284 142 287 144
rect 280 140 287 142
rect 218 133 223 138
rect 282 135 287 140
rect 289 135 294 146
rect 296 144 305 146
rect 333 145 339 147
rect 296 135 307 144
rect 309 142 316 144
rect 309 140 312 142
rect 314 140 316 142
rect 309 138 316 140
rect 322 143 329 145
rect 322 141 324 143
rect 326 141 329 143
rect 322 139 329 141
rect 331 143 339 145
rect 331 141 334 143
rect 336 141 339 143
rect 331 139 339 141
rect 341 139 346 147
rect 348 145 356 147
rect 348 143 351 145
rect 353 143 356 145
rect 348 139 356 143
rect 358 139 363 147
rect 365 145 373 147
rect 365 143 368 145
rect 370 143 373 145
rect 365 139 373 143
rect 309 135 314 138
rect 368 138 373 139
rect 375 144 380 147
rect 391 144 396 147
rect 375 142 382 144
rect 375 140 378 142
rect 380 140 382 142
rect 375 138 382 140
rect 389 142 396 144
rect 389 140 391 142
rect 393 140 396 142
rect 389 138 396 140
rect 398 145 406 147
rect 398 143 401 145
rect 403 143 406 145
rect 398 139 406 143
rect 408 139 413 147
rect 415 145 423 147
rect 415 143 418 145
rect 420 143 423 145
rect 415 139 423 143
rect 425 139 430 147
rect 432 145 438 147
rect 432 143 440 145
rect 432 141 435 143
rect 437 141 440 143
rect 432 139 440 141
rect 442 143 449 145
rect 458 144 463 147
rect 442 141 445 143
rect 447 141 449 143
rect 442 139 449 141
rect 456 142 463 144
rect 456 140 458 142
rect 460 140 463 142
rect 398 138 403 139
rect 456 138 463 140
rect 465 145 473 147
rect 465 143 468 145
rect 470 143 473 145
rect 465 139 473 143
rect 475 139 480 147
rect 482 145 490 147
rect 482 143 485 145
rect 487 143 490 145
rect 482 139 490 143
rect 492 139 497 147
rect 499 145 505 147
rect 564 154 570 156
rect 564 152 566 154
rect 568 152 570 154
rect 533 150 539 152
rect 533 148 535 150
rect 537 148 539 150
rect 499 143 507 145
rect 499 141 502 143
rect 504 141 507 143
rect 499 139 507 141
rect 509 143 516 145
rect 509 141 512 143
rect 514 141 516 143
rect 533 146 539 148
rect 552 150 558 152
rect 552 148 554 150
rect 556 148 558 150
rect 552 146 558 148
rect 533 142 537 146
rect 509 139 516 141
rect 524 139 529 142
rect 465 138 470 139
rect 522 137 529 139
rect 522 135 524 137
rect 526 135 529 137
rect 522 133 529 135
rect 531 139 537 142
rect 553 139 558 146
rect 531 133 539 139
rect 541 137 549 139
rect 541 135 544 137
rect 546 135 549 137
rect 541 133 549 135
rect 551 133 558 139
rect 564 150 570 152
rect 564 138 572 150
rect 574 138 579 150
rect 581 147 586 150
rect 581 144 589 147
rect 581 142 584 144
rect 586 142 589 144
rect 581 138 589 142
rect 591 142 599 147
rect 591 140 594 142
rect 596 140 599 142
rect 591 138 599 140
rect 601 145 610 147
rect 601 143 606 145
rect 608 143 610 145
rect 601 142 610 143
rect 601 138 615 142
rect 610 133 615 138
rect 617 139 622 142
rect 617 137 624 139
rect 617 135 620 137
rect 622 135 624 137
rect 617 133 624 135
rect 6 39 13 41
rect 6 37 8 39
rect 10 37 13 39
rect 6 35 13 37
rect 8 32 13 35
rect 15 35 23 41
rect 25 39 33 41
rect 25 37 28 39
rect 30 37 33 39
rect 25 35 33 37
rect 35 35 42 41
rect 95 39 102 41
rect 57 36 62 39
rect 15 32 21 35
rect 17 28 21 32
rect 37 28 42 35
rect 55 34 62 36
rect 55 32 57 34
rect 59 32 62 34
rect 55 30 62 32
rect 64 30 75 39
rect 17 26 23 28
rect 17 24 19 26
rect 21 24 23 26
rect 17 22 23 24
rect 36 26 42 28
rect 66 28 75 30
rect 77 28 82 39
rect 84 34 89 39
rect 95 37 97 39
rect 99 37 102 39
rect 95 35 102 37
rect 84 32 91 34
rect 97 32 102 35
rect 104 36 109 41
rect 209 39 216 41
rect 171 36 176 39
rect 104 32 118 36
rect 84 30 87 32
rect 89 30 91 32
rect 84 28 91 30
rect 109 31 118 32
rect 109 29 111 31
rect 113 29 118 31
rect 36 24 38 26
rect 40 24 42 26
rect 36 22 42 24
rect 66 22 73 28
rect 109 27 118 29
rect 120 34 128 36
rect 120 32 123 34
rect 125 32 128 34
rect 120 27 128 32
rect 130 32 138 36
rect 130 30 133 32
rect 135 30 138 32
rect 130 27 138 30
rect 66 20 68 22
rect 70 20 73 22
rect 66 18 73 20
rect 133 24 138 27
rect 140 24 145 36
rect 147 24 155 36
rect 169 34 176 36
rect 169 32 171 34
rect 173 32 176 34
rect 169 30 176 32
rect 178 30 189 39
rect 180 28 189 30
rect 191 28 196 39
rect 198 34 203 39
rect 209 37 211 39
rect 213 37 216 39
rect 209 35 216 37
rect 198 32 205 34
rect 211 32 216 35
rect 218 36 223 41
rect 218 32 232 36
rect 198 30 201 32
rect 203 30 205 32
rect 198 28 205 30
rect 223 31 232 32
rect 223 29 225 31
rect 227 29 232 31
rect 149 22 155 24
rect 149 20 151 22
rect 153 20 155 22
rect 149 18 155 20
rect 180 22 187 28
rect 223 27 232 29
rect 234 34 242 36
rect 234 32 237 34
rect 239 32 242 34
rect 234 27 242 32
rect 244 32 252 36
rect 244 30 247 32
rect 249 30 252 32
rect 244 27 252 30
rect 180 20 182 22
rect 184 20 187 22
rect 180 18 187 20
rect 247 24 252 27
rect 254 24 259 36
rect 261 24 269 36
rect 282 34 287 39
rect 280 32 287 34
rect 280 30 282 32
rect 284 30 287 32
rect 280 28 287 30
rect 289 28 294 39
rect 296 30 307 39
rect 309 36 314 39
rect 309 34 316 36
rect 368 35 373 36
rect 309 32 312 34
rect 314 32 316 34
rect 309 30 316 32
rect 322 33 329 35
rect 322 31 324 33
rect 326 31 329 33
rect 296 28 305 30
rect 263 22 269 24
rect 263 20 265 22
rect 267 20 269 22
rect 263 18 269 20
rect 298 22 305 28
rect 322 29 329 31
rect 331 33 339 35
rect 331 31 334 33
rect 336 31 339 33
rect 331 29 339 31
rect 298 20 301 22
rect 303 20 305 22
rect 298 18 305 20
rect 333 27 339 29
rect 341 27 346 35
rect 348 31 356 35
rect 348 29 351 31
rect 353 29 356 31
rect 348 27 356 29
rect 358 27 363 35
rect 365 31 373 35
rect 365 29 368 31
rect 370 29 373 31
rect 365 27 373 29
rect 375 34 382 36
rect 375 32 378 34
rect 380 32 382 34
rect 375 30 382 32
rect 389 34 396 36
rect 389 32 391 34
rect 393 32 396 34
rect 389 30 396 32
rect 375 27 380 30
rect 391 27 396 30
rect 398 35 403 36
rect 398 31 406 35
rect 398 29 401 31
rect 403 29 406 31
rect 398 27 406 29
rect 408 27 413 35
rect 415 31 423 35
rect 415 29 418 31
rect 420 29 423 31
rect 415 27 423 29
rect 425 27 430 35
rect 432 33 440 35
rect 432 31 435 33
rect 437 31 440 33
rect 432 29 440 31
rect 442 33 449 35
rect 442 31 445 33
rect 447 31 449 33
rect 442 29 449 31
rect 456 34 463 36
rect 456 32 458 34
rect 460 32 463 34
rect 456 30 463 32
rect 432 27 438 29
rect 458 27 463 30
rect 465 35 470 36
rect 522 39 529 41
rect 522 37 524 39
rect 526 37 529 39
rect 522 35 529 37
rect 465 31 473 35
rect 465 29 468 31
rect 470 29 473 31
rect 465 27 473 29
rect 475 27 480 35
rect 482 31 490 35
rect 482 29 485 31
rect 487 29 490 31
rect 482 27 490 29
rect 492 27 497 35
rect 499 33 507 35
rect 499 31 502 33
rect 504 31 507 33
rect 499 29 507 31
rect 509 33 516 35
rect 509 31 512 33
rect 514 31 516 33
rect 524 32 529 35
rect 531 35 539 41
rect 541 39 549 41
rect 541 37 544 39
rect 546 37 549 39
rect 541 35 549 37
rect 551 35 558 41
rect 610 36 615 41
rect 531 32 537 35
rect 509 29 516 31
rect 499 27 505 29
rect 533 28 537 32
rect 553 28 558 35
rect 533 26 539 28
rect 533 24 535 26
rect 537 24 539 26
rect 533 22 539 24
rect 552 26 558 28
rect 552 24 554 26
rect 556 24 558 26
rect 552 22 558 24
rect 564 24 572 36
rect 574 24 579 36
rect 581 32 589 36
rect 581 30 584 32
rect 586 30 589 32
rect 581 27 589 30
rect 591 34 599 36
rect 591 32 594 34
rect 596 32 599 34
rect 591 27 599 32
rect 601 32 615 36
rect 617 39 624 41
rect 617 37 620 39
rect 622 37 624 39
rect 617 35 624 37
rect 617 32 622 35
rect 601 31 610 32
rect 601 29 606 31
rect 608 29 610 31
rect 601 27 610 29
rect 581 24 586 27
rect 564 22 570 24
rect 564 20 566 22
rect 568 20 570 22
rect 564 18 570 20
<< pdif >>
rect 8 116 13 121
rect 6 114 13 116
rect 6 112 8 114
rect 10 112 13 114
rect 6 107 13 112
rect 6 105 8 107
rect 10 105 13 107
rect 6 103 13 105
rect 15 114 23 121
rect 55 118 62 120
rect 55 116 57 118
rect 59 116 62 118
rect 15 103 26 114
rect 17 97 26 103
rect 17 95 19 97
rect 21 95 26 97
rect 17 93 26 95
rect 28 93 33 114
rect 35 106 40 114
rect 55 111 62 116
rect 55 109 57 111
rect 59 109 62 111
rect 55 107 62 109
rect 35 104 42 106
rect 35 102 38 104
rect 40 102 42 104
rect 57 102 62 107
rect 64 113 70 120
rect 103 118 110 120
rect 103 116 105 118
rect 107 116 110 118
rect 103 114 110 116
rect 64 106 72 113
rect 64 104 67 106
rect 69 104 72 106
rect 64 102 72 104
rect 35 100 42 102
rect 35 93 40 100
rect 66 100 72 102
rect 74 111 82 113
rect 74 109 77 111
rect 79 109 82 111
rect 74 104 82 109
rect 74 102 77 104
rect 79 102 82 104
rect 74 100 82 102
rect 84 104 91 113
rect 84 102 87 104
rect 89 102 91 104
rect 84 100 91 102
rect 105 93 110 114
rect 112 104 126 120
rect 112 102 115 104
rect 117 102 126 104
rect 128 118 136 120
rect 128 116 131 118
rect 133 116 136 118
rect 128 111 136 116
rect 128 109 131 111
rect 133 109 136 111
rect 128 102 136 109
rect 138 111 146 120
rect 138 109 141 111
rect 143 109 146 111
rect 138 102 146 109
rect 112 97 124 102
rect 112 95 115 97
rect 117 95 124 97
rect 112 93 124 95
rect 141 93 146 102
rect 148 105 153 120
rect 169 118 176 120
rect 169 116 171 118
rect 173 116 176 118
rect 169 111 176 116
rect 169 109 171 111
rect 173 109 176 111
rect 169 107 176 109
rect 148 103 155 105
rect 148 101 151 103
rect 153 101 155 103
rect 171 102 176 107
rect 178 113 184 120
rect 217 118 224 120
rect 217 116 219 118
rect 221 116 224 118
rect 217 114 224 116
rect 178 106 186 113
rect 178 104 181 106
rect 183 104 186 106
rect 178 102 186 104
rect 148 99 155 101
rect 148 93 153 99
rect 180 100 186 102
rect 188 111 196 113
rect 188 109 191 111
rect 193 109 196 111
rect 188 104 196 109
rect 188 102 191 104
rect 193 102 196 104
rect 188 100 196 102
rect 198 104 205 113
rect 198 102 201 104
rect 203 102 205 104
rect 198 100 205 102
rect 219 93 224 114
rect 226 104 240 120
rect 226 102 229 104
rect 231 102 240 104
rect 242 118 250 120
rect 242 116 245 118
rect 247 116 250 118
rect 242 111 250 116
rect 242 109 245 111
rect 247 109 250 111
rect 242 102 250 109
rect 252 111 260 120
rect 252 109 255 111
rect 257 109 260 111
rect 252 102 260 109
rect 226 97 238 102
rect 226 95 229 97
rect 231 95 238 97
rect 226 93 238 95
rect 255 93 260 102
rect 262 105 267 120
rect 301 113 307 120
rect 262 103 269 105
rect 262 101 265 103
rect 267 101 269 103
rect 262 99 269 101
rect 280 104 287 113
rect 280 102 282 104
rect 284 102 287 104
rect 280 100 287 102
rect 289 111 297 113
rect 289 109 292 111
rect 294 109 297 111
rect 289 104 297 109
rect 289 102 292 104
rect 294 102 297 104
rect 289 100 297 102
rect 299 106 307 113
rect 299 104 302 106
rect 304 104 307 106
rect 299 102 307 104
rect 309 118 316 120
rect 309 116 312 118
rect 314 116 316 118
rect 309 111 316 116
rect 322 119 329 121
rect 322 117 324 119
rect 326 117 329 119
rect 322 115 329 117
rect 324 113 329 115
rect 331 113 337 121
rect 309 109 312 111
rect 314 109 316 111
rect 309 107 316 109
rect 333 109 337 113
rect 368 109 373 111
rect 309 102 314 107
rect 333 105 339 109
rect 299 100 305 102
rect 262 93 267 99
rect 332 97 339 105
rect 332 95 334 97
rect 336 95 339 97
rect 332 93 339 95
rect 341 93 346 109
rect 348 107 356 109
rect 348 105 351 107
rect 353 105 356 107
rect 348 93 356 105
rect 358 93 363 109
rect 365 97 373 109
rect 365 95 368 97
rect 370 95 373 97
rect 365 93 373 95
rect 375 106 380 111
rect 391 106 396 111
rect 375 104 382 106
rect 375 102 378 104
rect 380 102 382 104
rect 375 100 382 102
rect 389 104 396 106
rect 389 102 391 104
rect 393 102 396 104
rect 389 100 396 102
rect 375 93 380 100
rect 391 93 396 100
rect 398 109 403 111
rect 434 113 440 121
rect 442 119 449 121
rect 442 117 445 119
rect 447 117 449 119
rect 442 115 449 117
rect 442 113 447 115
rect 434 109 438 113
rect 398 97 406 109
rect 398 95 401 97
rect 403 95 406 97
rect 398 93 406 95
rect 408 93 413 109
rect 415 107 423 109
rect 415 105 418 107
rect 420 105 423 107
rect 415 93 423 105
rect 425 93 430 109
rect 432 105 438 109
rect 458 106 463 111
rect 432 97 439 105
rect 456 104 463 106
rect 456 102 458 104
rect 460 102 463 104
rect 456 100 463 102
rect 432 95 435 97
rect 437 95 439 97
rect 432 93 439 95
rect 458 93 463 100
rect 465 109 470 111
rect 501 113 507 121
rect 509 119 516 121
rect 509 117 512 119
rect 514 117 516 119
rect 509 115 516 117
rect 524 116 529 121
rect 509 113 514 115
rect 522 114 529 116
rect 501 109 505 113
rect 465 97 473 109
rect 465 95 468 97
rect 470 95 473 97
rect 465 93 473 95
rect 475 93 480 109
rect 482 107 490 109
rect 482 105 485 107
rect 487 105 490 107
rect 482 93 490 105
rect 492 93 497 109
rect 499 105 505 109
rect 522 112 524 114
rect 526 112 529 114
rect 499 97 506 105
rect 522 107 529 112
rect 522 105 524 107
rect 526 105 529 107
rect 522 103 529 105
rect 531 114 539 121
rect 531 103 542 114
rect 499 95 502 97
rect 504 95 506 97
rect 533 97 542 103
rect 499 93 506 95
rect 533 95 535 97
rect 537 95 542 97
rect 533 93 542 95
rect 544 93 549 114
rect 551 106 556 114
rect 551 104 558 106
rect 566 105 571 120
rect 551 102 554 104
rect 556 102 558 104
rect 551 100 558 102
rect 564 103 571 105
rect 564 101 566 103
rect 568 101 571 103
rect 551 93 556 100
rect 564 99 571 101
rect 566 93 571 99
rect 573 111 581 120
rect 573 109 576 111
rect 578 109 581 111
rect 573 102 581 109
rect 583 118 591 120
rect 583 116 586 118
rect 588 116 591 118
rect 583 111 591 116
rect 583 109 586 111
rect 588 109 591 111
rect 583 102 591 109
rect 593 104 607 120
rect 593 102 602 104
rect 604 102 607 104
rect 573 93 578 102
rect 595 97 607 102
rect 595 95 602 97
rect 604 95 607 97
rect 595 93 607 95
rect 609 118 616 120
rect 609 116 612 118
rect 614 116 616 118
rect 609 114 616 116
rect 609 93 614 114
rect 17 79 26 81
rect 17 77 19 79
rect 21 77 26 79
rect 17 71 26 77
rect 6 69 13 71
rect 6 67 8 69
rect 10 67 13 69
rect 6 62 13 67
rect 6 60 8 62
rect 10 60 13 62
rect 6 58 13 60
rect 8 53 13 58
rect 15 60 26 71
rect 28 60 33 81
rect 35 74 40 81
rect 35 72 42 74
rect 66 72 72 74
rect 35 70 38 72
rect 40 70 42 72
rect 35 68 42 70
rect 35 60 40 68
rect 57 67 62 72
rect 55 65 62 67
rect 55 63 57 65
rect 59 63 62 65
rect 15 53 23 60
rect 55 58 62 63
rect 55 56 57 58
rect 59 56 62 58
rect 55 54 62 56
rect 64 70 72 72
rect 64 68 67 70
rect 69 68 72 70
rect 64 61 72 68
rect 74 72 82 74
rect 74 70 77 72
rect 79 70 82 72
rect 74 65 82 70
rect 74 63 77 65
rect 79 63 82 65
rect 74 61 82 63
rect 84 72 91 74
rect 84 70 87 72
rect 89 70 91 72
rect 84 61 91 70
rect 64 54 70 61
rect 105 60 110 81
rect 103 58 110 60
rect 103 56 105 58
rect 107 56 110 58
rect 103 54 110 56
rect 112 79 124 81
rect 112 77 115 79
rect 117 77 124 79
rect 112 72 124 77
rect 141 72 146 81
rect 112 70 115 72
rect 117 70 126 72
rect 112 54 126 70
rect 128 65 136 72
rect 128 63 131 65
rect 133 63 136 65
rect 128 58 136 63
rect 128 56 131 58
rect 133 56 136 58
rect 128 54 136 56
rect 138 65 146 72
rect 138 63 141 65
rect 143 63 146 65
rect 138 54 146 63
rect 148 75 153 81
rect 148 73 155 75
rect 148 71 151 73
rect 153 71 155 73
rect 180 72 186 74
rect 148 69 155 71
rect 148 54 153 69
rect 171 67 176 72
rect 169 65 176 67
rect 169 63 171 65
rect 173 63 176 65
rect 169 58 176 63
rect 169 56 171 58
rect 173 56 176 58
rect 169 54 176 56
rect 178 70 186 72
rect 178 68 181 70
rect 183 68 186 70
rect 178 61 186 68
rect 188 72 196 74
rect 188 70 191 72
rect 193 70 196 72
rect 188 65 196 70
rect 188 63 191 65
rect 193 63 196 65
rect 188 61 196 63
rect 198 72 205 74
rect 198 70 201 72
rect 203 70 205 72
rect 198 61 205 70
rect 178 54 184 61
rect 219 60 224 81
rect 217 58 224 60
rect 217 56 219 58
rect 221 56 224 58
rect 217 54 224 56
rect 226 79 238 81
rect 226 77 229 79
rect 231 77 238 79
rect 226 72 238 77
rect 255 72 260 81
rect 226 70 229 72
rect 231 70 240 72
rect 226 54 240 70
rect 242 65 250 72
rect 242 63 245 65
rect 247 63 250 65
rect 242 58 250 63
rect 242 56 245 58
rect 247 56 250 58
rect 242 54 250 56
rect 252 65 260 72
rect 252 63 255 65
rect 257 63 260 65
rect 252 54 260 63
rect 262 75 267 81
rect 262 73 269 75
rect 332 79 339 81
rect 332 77 334 79
rect 336 77 339 79
rect 262 71 265 73
rect 267 71 269 73
rect 262 69 269 71
rect 280 72 287 74
rect 280 70 282 72
rect 284 70 287 72
rect 262 54 267 69
rect 280 61 287 70
rect 289 72 297 74
rect 289 70 292 72
rect 294 70 297 72
rect 289 65 297 70
rect 289 63 292 65
rect 294 63 297 65
rect 289 61 297 63
rect 299 72 305 74
rect 299 70 307 72
rect 299 68 302 70
rect 304 68 307 70
rect 299 61 307 68
rect 301 54 307 61
rect 309 67 314 72
rect 332 69 339 77
rect 309 65 316 67
rect 309 63 312 65
rect 314 63 316 65
rect 309 58 316 63
rect 333 65 339 69
rect 341 65 346 81
rect 348 69 356 81
rect 348 67 351 69
rect 353 67 356 69
rect 348 65 356 67
rect 358 65 363 81
rect 365 79 373 81
rect 365 77 368 79
rect 370 77 373 79
rect 365 65 373 77
rect 333 61 337 65
rect 324 59 329 61
rect 309 56 312 58
rect 314 56 316 58
rect 309 54 316 56
rect 322 57 329 59
rect 322 55 324 57
rect 326 55 329 57
rect 322 53 329 55
rect 331 53 337 61
rect 368 63 373 65
rect 375 74 380 81
rect 391 74 396 81
rect 375 72 382 74
rect 375 70 378 72
rect 380 70 382 72
rect 375 68 382 70
rect 389 72 396 74
rect 389 70 391 72
rect 393 70 396 72
rect 389 68 396 70
rect 375 63 380 68
rect 391 63 396 68
rect 398 79 406 81
rect 398 77 401 79
rect 403 77 406 79
rect 398 65 406 77
rect 408 65 413 81
rect 415 69 423 81
rect 415 67 418 69
rect 420 67 423 69
rect 415 65 423 67
rect 425 65 430 81
rect 432 79 439 81
rect 432 77 435 79
rect 437 77 439 79
rect 432 69 439 77
rect 458 74 463 81
rect 456 72 463 74
rect 456 70 458 72
rect 460 70 463 72
rect 432 65 438 69
rect 456 68 463 70
rect 398 63 403 65
rect 434 61 438 65
rect 458 63 463 68
rect 465 79 473 81
rect 465 77 468 79
rect 470 77 473 79
rect 465 65 473 77
rect 475 65 480 81
rect 482 69 490 81
rect 482 67 485 69
rect 487 67 490 69
rect 482 65 490 67
rect 492 65 497 81
rect 499 79 506 81
rect 499 77 502 79
rect 504 77 506 79
rect 533 79 542 81
rect 499 69 506 77
rect 533 77 535 79
rect 537 77 542 79
rect 533 71 542 77
rect 499 65 505 69
rect 465 63 470 65
rect 434 53 440 61
rect 442 59 447 61
rect 442 57 449 59
rect 442 55 445 57
rect 447 55 449 57
rect 442 53 449 55
rect 501 61 505 65
rect 522 69 529 71
rect 522 67 524 69
rect 526 67 529 69
rect 522 62 529 67
rect 501 53 507 61
rect 509 59 514 61
rect 522 60 524 62
rect 526 60 529 62
rect 509 57 516 59
rect 522 58 529 60
rect 509 55 512 57
rect 514 55 516 57
rect 509 53 516 55
rect 524 53 529 58
rect 531 60 542 71
rect 544 60 549 81
rect 551 74 556 81
rect 566 75 571 81
rect 551 72 558 74
rect 551 70 554 72
rect 556 70 558 72
rect 551 68 558 70
rect 564 73 571 75
rect 564 71 566 73
rect 568 71 571 73
rect 564 69 571 71
rect 551 60 556 68
rect 531 53 539 60
rect 566 54 571 69
rect 573 72 578 81
rect 595 79 607 81
rect 595 77 602 79
rect 604 77 607 79
rect 595 72 607 77
rect 573 65 581 72
rect 573 63 576 65
rect 578 63 581 65
rect 573 54 581 63
rect 583 65 591 72
rect 583 63 586 65
rect 588 63 591 65
rect 583 58 591 63
rect 583 56 586 58
rect 588 56 591 58
rect 583 54 591 56
rect 593 70 602 72
rect 604 70 607 72
rect 593 54 607 70
rect 609 60 614 81
rect 609 58 616 60
rect 609 56 612 58
rect 614 56 616 58
rect 609 54 616 56
<< alu1 >>
rect 2 154 632 159
rect 2 152 9 154
rect 11 152 58 154
rect 60 152 68 154
rect 70 152 98 154
rect 100 152 151 154
rect 153 152 172 154
rect 174 152 182 154
rect 184 152 212 154
rect 214 152 265 154
rect 267 152 301 154
rect 303 152 311 154
rect 313 152 525 154
rect 527 152 566 154
rect 568 152 619 154
rect 621 152 632 154
rect 2 151 632 152
rect 55 142 67 146
rect 55 140 57 142
rect 59 140 67 142
rect 131 144 155 145
rect 6 137 11 139
rect 6 135 8 137
rect 10 135 11 137
rect 6 133 11 135
rect 6 114 10 133
rect 38 129 42 138
rect 6 112 8 114
rect 6 107 10 112
rect 6 105 8 107
rect 21 128 42 129
rect 21 126 25 128
rect 27 126 39 128
rect 41 126 42 128
rect 21 125 42 126
rect 21 119 35 121
rect 37 119 42 121
rect 21 117 42 119
rect 38 115 42 117
rect 55 120 59 140
rect 131 142 133 144
rect 135 142 155 144
rect 131 141 155 142
rect 79 137 84 138
rect 79 135 80 137
rect 82 135 84 137
rect 79 129 84 135
rect 55 118 60 120
rect 55 116 57 118
rect 59 116 60 118
rect 55 115 60 116
rect 38 111 60 115
rect 38 108 42 111
rect 55 109 57 111
rect 59 109 60 111
rect 70 128 84 129
rect 70 126 74 128
rect 76 126 84 128
rect 70 125 84 126
rect 103 137 116 138
rect 103 135 105 137
rect 107 135 116 137
rect 103 133 116 135
rect 103 132 113 133
rect 111 131 113 132
rect 115 131 116 133
rect 78 120 91 121
rect 78 118 84 120
rect 86 118 91 120
rect 78 117 91 118
rect 55 107 60 109
rect 6 101 19 105
rect 6 100 10 101
rect 87 113 91 117
rect 87 111 88 113
rect 90 111 91 113
rect 87 108 91 111
rect 95 120 100 122
rect 95 118 97 120
rect 99 118 100 120
rect 95 113 100 118
rect 111 124 116 131
rect 151 136 155 141
rect 151 134 152 136
rect 154 134 155 136
rect 95 111 97 113
rect 99 111 100 113
rect 95 106 100 111
rect 95 100 107 106
rect 151 113 155 134
rect 139 111 155 113
rect 139 109 141 111
rect 143 109 155 111
rect 139 108 155 109
rect 169 142 181 146
rect 169 140 171 142
rect 173 140 181 142
rect 245 144 269 145
rect 169 128 173 140
rect 245 142 247 144
rect 249 142 269 144
rect 245 141 269 142
rect 169 126 170 128
rect 172 126 173 128
rect 169 120 173 126
rect 193 137 198 138
rect 193 135 194 137
rect 196 135 198 137
rect 193 129 198 135
rect 169 118 174 120
rect 169 116 171 118
rect 173 116 174 118
rect 169 111 174 116
rect 169 109 171 111
rect 173 109 174 111
rect 184 128 198 129
rect 184 126 188 128
rect 190 126 198 128
rect 184 125 198 126
rect 217 137 230 138
rect 217 135 219 137
rect 221 135 230 137
rect 217 133 230 135
rect 217 132 227 133
rect 225 131 227 132
rect 229 131 230 133
rect 192 120 205 121
rect 192 118 198 120
rect 200 118 205 120
rect 192 117 205 118
rect 201 114 205 117
rect 209 120 214 122
rect 209 118 211 120
rect 213 118 214 120
rect 209 114 214 118
rect 225 124 230 131
rect 169 107 174 109
rect 201 113 214 114
rect 201 111 202 113
rect 204 111 211 113
rect 213 111 214 113
rect 201 110 214 111
rect 201 108 205 110
rect 209 106 214 110
rect 209 104 221 106
rect 209 102 211 104
rect 213 102 221 104
rect 209 100 221 102
rect 201 95 205 100
rect 265 121 269 141
rect 287 129 292 138
rect 304 142 316 146
rect 304 140 312 142
rect 314 140 316 142
rect 287 128 301 129
rect 287 126 295 128
rect 297 126 301 128
rect 287 125 301 126
rect 265 119 266 121
rect 268 119 269 121
rect 265 113 269 119
rect 253 111 269 113
rect 253 109 255 111
rect 257 109 269 111
rect 253 108 269 109
rect 280 120 293 121
rect 280 118 285 120
rect 287 118 293 120
rect 280 117 293 118
rect 280 108 284 117
rect 312 136 316 140
rect 312 134 313 136
rect 315 134 316 136
rect 312 120 316 134
rect 311 118 316 120
rect 311 116 312 118
rect 314 116 316 118
rect 378 144 382 146
rect 377 142 382 144
rect 377 140 378 142
rect 380 140 382 142
rect 377 138 382 140
rect 329 136 342 137
rect 329 134 330 136
rect 332 134 342 136
rect 329 133 342 134
rect 336 128 342 133
rect 336 126 337 128
rect 339 126 342 128
rect 336 124 342 126
rect 362 123 366 130
rect 362 122 364 123
rect 354 121 364 122
rect 354 120 366 121
rect 354 118 355 120
rect 357 118 366 120
rect 354 116 366 118
rect 311 111 316 116
rect 311 109 312 111
rect 314 109 316 111
rect 311 107 316 109
rect 322 112 335 113
rect 322 110 332 112
rect 334 110 335 112
rect 322 109 335 110
rect 322 108 327 109
rect 378 128 382 138
rect 378 126 379 128
rect 381 126 382 128
rect 322 106 324 108
rect 326 106 327 108
rect 322 100 327 106
rect 378 105 382 126
rect 369 104 382 105
rect 369 102 378 104
rect 380 102 382 104
rect 369 101 382 102
rect 389 144 393 146
rect 389 142 394 144
rect 389 140 391 142
rect 393 140 394 142
rect 456 144 460 146
rect 389 138 394 140
rect 389 105 393 138
rect 429 136 442 137
rect 405 128 409 130
rect 405 126 406 128
rect 408 126 409 128
rect 405 123 409 126
rect 407 122 409 123
rect 407 121 417 122
rect 405 116 417 121
rect 429 134 437 136
rect 439 134 442 136
rect 429 133 442 134
rect 429 128 435 133
rect 429 126 432 128
rect 434 126 435 128
rect 429 124 435 126
rect 456 142 461 144
rect 456 140 458 142
rect 460 140 461 142
rect 564 144 588 145
rect 456 138 461 140
rect 456 136 460 138
rect 456 134 457 136
rect 459 134 460 136
rect 496 136 509 137
rect 436 109 449 113
rect 444 108 449 109
rect 389 104 402 105
rect 444 106 445 108
rect 447 106 449 108
rect 389 102 391 104
rect 393 102 402 104
rect 389 101 402 102
rect 444 100 449 106
rect 456 105 460 134
rect 472 123 476 130
rect 474 122 476 123
rect 474 121 484 122
rect 472 119 480 121
rect 482 119 484 121
rect 472 116 484 119
rect 496 134 505 136
rect 507 134 509 136
rect 496 133 509 134
rect 496 128 502 133
rect 496 126 499 128
rect 501 126 502 128
rect 496 124 502 126
rect 564 142 584 144
rect 586 142 588 144
rect 564 141 588 142
rect 522 137 527 139
rect 522 135 524 137
rect 526 135 527 137
rect 522 133 527 135
rect 522 120 526 133
rect 522 118 523 120
rect 525 118 526 120
rect 522 114 526 118
rect 554 129 558 138
rect 503 112 516 113
rect 503 110 504 112
rect 506 110 516 112
rect 503 109 516 110
rect 511 108 516 109
rect 456 104 469 105
rect 511 106 512 108
rect 514 106 516 108
rect 456 102 458 104
rect 460 102 469 104
rect 456 101 469 102
rect 511 100 516 106
rect 522 112 524 114
rect 522 107 526 112
rect 522 105 524 107
rect 537 128 558 129
rect 537 126 541 128
rect 543 126 558 128
rect 537 125 558 126
rect 564 136 568 141
rect 564 134 565 136
rect 567 134 568 136
rect 537 119 551 121
rect 553 119 558 121
rect 537 117 558 119
rect 554 108 558 117
rect 564 113 568 134
rect 603 133 616 138
rect 603 131 604 133
rect 606 132 616 133
rect 606 131 608 132
rect 564 111 580 113
rect 564 109 576 111
rect 578 109 580 111
rect 564 108 580 109
rect 603 124 608 131
rect 619 120 624 122
rect 619 118 620 120
rect 622 118 624 120
rect 522 101 535 105
rect 619 106 624 118
rect 522 100 526 101
rect 612 100 624 106
rect 2 94 632 95
rect 2 92 9 94
rect 11 92 58 94
rect 60 92 131 94
rect 133 92 172 94
rect 174 92 245 94
rect 247 92 311 94
rect 313 92 525 94
rect 527 92 586 94
rect 588 92 632 94
rect 2 82 632 92
rect 2 80 9 82
rect 11 80 58 82
rect 60 80 131 82
rect 133 80 172 82
rect 174 80 245 82
rect 247 80 311 82
rect 313 80 525 82
rect 527 80 586 82
rect 588 80 632 82
rect 2 79 632 80
rect 6 73 10 74
rect 6 69 19 73
rect 6 67 8 69
rect 6 62 10 67
rect 6 60 8 62
rect 6 57 10 60
rect 38 63 42 66
rect 55 65 60 67
rect 55 63 57 65
rect 59 63 60 65
rect 95 68 107 74
rect 6 55 7 57
rect 9 55 10 57
rect 6 41 10 55
rect 38 59 60 63
rect 38 57 42 59
rect 21 55 42 57
rect 21 53 35 55
rect 37 53 42 55
rect 55 58 60 59
rect 55 56 57 58
rect 59 56 60 58
rect 55 54 60 56
rect 87 63 91 66
rect 87 61 88 63
rect 90 61 91 63
rect 6 39 11 41
rect 6 37 8 39
rect 10 37 11 39
rect 6 35 11 37
rect 21 48 42 49
rect 21 46 25 48
rect 27 46 39 48
rect 41 46 42 48
rect 21 45 42 46
rect 38 36 42 45
rect 55 34 59 54
rect 87 57 91 61
rect 78 56 91 57
rect 78 54 84 56
rect 86 54 91 56
rect 78 53 91 54
rect 95 63 100 68
rect 95 61 97 63
rect 99 61 100 63
rect 95 56 100 61
rect 95 54 97 56
rect 99 54 100 56
rect 95 52 100 54
rect 70 48 84 49
rect 70 46 74 48
rect 76 46 84 48
rect 70 45 84 46
rect 55 32 57 34
rect 59 32 67 34
rect 55 28 67 32
rect 79 39 84 45
rect 79 37 80 39
rect 82 37 84 39
rect 79 36 84 37
rect 111 43 116 50
rect 139 65 155 66
rect 139 63 141 65
rect 143 63 155 65
rect 139 61 155 63
rect 111 42 113 43
rect 103 41 113 42
rect 115 41 116 43
rect 103 39 116 41
rect 103 37 105 39
rect 107 37 116 39
rect 103 36 116 37
rect 151 40 155 61
rect 151 38 152 40
rect 154 38 155 40
rect 151 33 155 38
rect 131 32 155 33
rect 131 30 133 32
rect 135 30 155 32
rect 131 29 155 30
rect 169 65 174 67
rect 169 63 171 65
rect 173 63 174 65
rect 209 68 221 74
rect 169 58 174 63
rect 169 56 171 58
rect 173 56 174 58
rect 169 54 174 56
rect 201 63 205 66
rect 201 61 202 63
rect 204 61 205 63
rect 169 48 173 54
rect 169 46 170 48
rect 172 46 173 48
rect 169 34 173 46
rect 201 57 205 61
rect 192 56 205 57
rect 192 54 198 56
rect 200 54 205 56
rect 192 53 205 54
rect 209 63 214 68
rect 209 61 211 63
rect 213 61 214 63
rect 209 56 214 61
rect 209 54 211 56
rect 213 54 214 56
rect 209 52 214 54
rect 184 48 198 49
rect 184 46 188 48
rect 190 46 198 48
rect 184 45 198 46
rect 169 32 171 34
rect 173 32 181 34
rect 169 28 181 32
rect 193 39 198 45
rect 193 37 194 39
rect 196 37 198 39
rect 193 36 198 37
rect 225 43 230 50
rect 253 65 269 66
rect 253 63 255 65
rect 257 63 269 65
rect 253 61 269 63
rect 265 55 269 61
rect 265 53 266 55
rect 268 53 269 55
rect 280 57 284 66
rect 322 68 327 74
rect 369 72 382 73
rect 369 70 378 72
rect 380 70 382 72
rect 311 65 316 67
rect 280 56 293 57
rect 280 54 285 56
rect 287 54 293 56
rect 280 53 293 54
rect 225 42 227 43
rect 217 41 227 42
rect 229 41 230 43
rect 217 39 230 41
rect 217 37 219 39
rect 221 37 230 39
rect 217 36 230 37
rect 265 33 269 53
rect 287 48 301 49
rect 287 46 295 48
rect 297 46 301 48
rect 287 45 301 46
rect 311 63 312 65
rect 314 63 316 65
rect 311 58 316 63
rect 322 66 324 68
rect 326 66 327 68
rect 369 69 382 70
rect 322 65 327 66
rect 322 64 335 65
rect 322 62 332 64
rect 334 62 335 64
rect 322 61 335 62
rect 311 56 312 58
rect 314 56 316 58
rect 311 54 316 56
rect 287 36 292 45
rect 312 40 316 54
rect 312 38 313 40
rect 315 38 316 40
rect 312 34 316 38
rect 245 32 269 33
rect 245 30 247 32
rect 249 30 269 32
rect 245 29 269 30
rect 304 32 312 34
rect 314 32 316 34
rect 304 28 316 32
rect 336 48 342 50
rect 336 46 337 48
rect 339 46 342 48
rect 336 41 342 46
rect 329 40 342 41
rect 329 38 330 40
rect 332 38 342 40
rect 354 56 366 58
rect 354 54 355 56
rect 357 54 366 56
rect 354 53 366 54
rect 354 52 364 53
rect 362 51 364 52
rect 362 44 366 51
rect 378 48 382 69
rect 378 46 379 48
rect 381 46 382 48
rect 329 37 342 38
rect 378 36 382 46
rect 377 34 382 36
rect 377 32 378 34
rect 380 32 382 34
rect 377 30 382 32
rect 378 28 382 30
rect 389 72 402 73
rect 389 70 391 72
rect 393 70 402 72
rect 389 69 402 70
rect 389 36 393 69
rect 444 68 449 74
rect 444 66 445 68
rect 447 66 449 68
rect 444 65 449 66
rect 436 61 449 65
rect 456 72 469 73
rect 456 70 458 72
rect 460 70 469 72
rect 456 69 469 70
rect 405 53 417 58
rect 407 52 417 53
rect 407 51 409 52
rect 405 48 409 51
rect 405 46 406 48
rect 408 46 409 48
rect 405 44 409 46
rect 429 48 435 50
rect 429 46 432 48
rect 434 46 435 48
rect 429 41 435 46
rect 429 40 442 41
rect 429 38 437 40
rect 439 38 442 40
rect 429 37 442 38
rect 389 34 394 36
rect 389 32 391 34
rect 393 32 394 34
rect 389 30 394 32
rect 389 28 393 30
rect 456 40 460 69
rect 511 68 516 74
rect 511 66 512 68
rect 514 66 516 68
rect 511 65 516 66
rect 503 64 516 65
rect 503 62 504 64
rect 506 62 516 64
rect 503 61 516 62
rect 522 73 526 74
rect 522 69 535 73
rect 522 67 524 69
rect 522 62 526 67
rect 522 60 524 62
rect 472 55 484 58
rect 472 53 480 55
rect 482 53 484 55
rect 474 52 484 53
rect 474 51 476 52
rect 456 38 457 40
rect 459 38 460 40
rect 472 44 476 51
rect 456 36 460 38
rect 496 48 502 50
rect 496 46 499 48
rect 501 46 502 48
rect 496 41 502 46
rect 496 40 509 41
rect 496 38 505 40
rect 507 38 509 40
rect 496 37 509 38
rect 456 34 461 36
rect 456 32 458 34
rect 460 32 461 34
rect 456 30 461 32
rect 456 28 460 30
rect 522 56 526 60
rect 522 54 523 56
rect 525 54 526 56
rect 522 41 526 54
rect 554 57 558 66
rect 537 55 558 57
rect 537 53 551 55
rect 553 53 558 55
rect 564 65 580 66
rect 564 63 576 65
rect 578 63 580 65
rect 564 61 580 63
rect 522 39 527 41
rect 522 37 524 39
rect 526 37 527 39
rect 522 35 527 37
rect 537 48 558 49
rect 537 46 541 48
rect 543 46 558 48
rect 537 45 558 46
rect 554 36 558 45
rect 564 40 568 61
rect 612 68 624 74
rect 564 38 565 40
rect 567 38 568 40
rect 564 33 568 38
rect 603 43 608 50
rect 619 56 624 68
rect 619 54 620 56
rect 622 54 624 56
rect 619 52 624 54
rect 603 41 604 43
rect 606 42 608 43
rect 606 41 616 42
rect 603 36 616 41
rect 564 32 588 33
rect 564 30 584 32
rect 586 30 588 32
rect 564 29 588 30
rect 2 22 632 23
rect 2 20 9 22
rect 11 20 58 22
rect 60 20 68 22
rect 70 20 98 22
rect 100 20 151 22
rect 153 20 172 22
rect 174 20 182 22
rect 184 20 212 22
rect 214 20 265 22
rect 267 20 301 22
rect 303 20 311 22
rect 313 20 525 22
rect 527 20 566 22
rect 568 20 619 22
rect 621 20 632 22
rect 2 15 632 20
<< alu2 >>
rect 79 137 111 138
rect 79 135 80 137
rect 82 135 105 137
rect 107 135 111 137
rect 79 133 111 135
rect 151 137 225 138
rect 151 136 194 137
rect 151 134 152 136
rect 154 135 194 136
rect 196 135 219 137
rect 221 135 225 137
rect 154 134 225 135
rect 151 133 225 134
rect 312 136 333 137
rect 312 134 313 136
rect 315 134 330 136
rect 332 134 333 136
rect 312 133 333 134
rect 436 136 460 137
rect 436 134 437 136
rect 439 134 457 136
rect 459 134 460 136
rect 436 133 460 134
rect 504 136 568 137
rect 504 134 505 136
rect 507 134 565 136
rect 567 134 568 136
rect 504 133 568 134
rect 38 128 173 129
rect 38 126 39 128
rect 41 126 170 128
rect 172 126 173 128
rect 38 125 173 126
rect 378 128 409 129
rect 378 126 379 128
rect 381 126 406 128
rect 408 126 409 128
rect 378 125 409 126
rect 265 121 359 122
rect 265 119 266 121
rect 268 120 359 121
rect 268 119 355 120
rect 265 118 355 119
rect 357 118 359 120
rect 265 117 359 118
rect 479 121 526 122
rect 479 119 480 121
rect 482 120 526 121
rect 482 119 523 120
rect 479 118 523 119
rect 525 118 526 120
rect 479 117 526 118
rect 87 113 100 114
rect 87 111 88 113
rect 90 111 97 113
rect 99 111 100 113
rect 87 110 100 111
rect 201 113 214 114
rect 201 111 202 113
rect 204 111 211 113
rect 213 111 214 113
rect 201 110 214 111
rect 331 112 508 113
rect 331 110 332 112
rect 334 110 504 112
rect 506 110 508 112
rect 201 100 205 110
rect 331 109 508 110
rect 210 104 214 105
rect 210 102 211 104
rect 213 102 214 104
rect 6 83 10 87
rect 210 83 214 102
rect 6 79 214 83
rect 6 57 10 79
rect 331 64 508 65
rect 87 63 100 64
rect 87 61 88 63
rect 90 61 97 63
rect 99 61 100 63
rect 87 60 100 61
rect 201 63 214 64
rect 201 61 202 63
rect 204 61 211 63
rect 213 61 214 63
rect 331 62 332 64
rect 334 62 504 64
rect 506 62 508 64
rect 331 61 508 62
rect 201 60 214 61
rect 6 55 7 57
rect 9 55 10 57
rect 6 54 10 55
rect 265 56 359 57
rect 265 55 355 56
rect 265 53 266 55
rect 268 54 355 55
rect 357 54 359 56
rect 268 53 359 54
rect 265 52 359 53
rect 479 56 526 57
rect 479 55 523 56
rect 479 53 480 55
rect 482 54 523 55
rect 525 54 526 56
rect 482 53 526 54
rect 479 52 526 53
rect 38 48 173 49
rect 38 46 39 48
rect 41 46 170 48
rect 172 46 173 48
rect 38 45 173 46
rect 378 48 409 49
rect 378 46 379 48
rect 381 46 406 48
rect 408 46 409 48
rect 378 45 409 46
rect 79 39 111 41
rect 79 37 80 39
rect 82 37 105 39
rect 107 37 111 39
rect 79 36 111 37
rect 151 40 225 41
rect 151 38 152 40
rect 154 39 225 40
rect 154 38 194 39
rect 151 37 194 38
rect 196 37 219 39
rect 221 37 225 39
rect 312 40 333 41
rect 312 38 313 40
rect 315 38 330 40
rect 332 38 333 40
rect 312 37 333 38
rect 436 40 460 41
rect 436 38 437 40
rect 439 38 457 40
rect 459 38 460 40
rect 436 37 460 38
rect 504 40 568 41
rect 504 38 505 40
rect 507 38 565 40
rect 567 38 568 40
rect 504 37 568 38
rect 151 36 225 37
<< ptie >>
rect 7 154 13 156
rect 7 152 9 154
rect 11 152 13 154
rect 56 154 62 156
rect 56 152 58 154
rect 60 152 62 154
rect 7 150 13 152
rect 56 150 62 152
rect 96 154 102 156
rect 96 152 98 154
rect 100 152 102 154
rect 96 150 102 152
rect 170 154 176 156
rect 170 152 172 154
rect 174 152 176 154
rect 170 150 176 152
rect 210 154 216 156
rect 210 152 212 154
rect 214 152 216 154
rect 210 150 216 152
rect 309 154 315 156
rect 309 152 311 154
rect 313 152 315 154
rect 309 150 315 152
rect 523 154 529 156
rect 523 152 525 154
rect 527 152 529 154
rect 523 150 529 152
rect 617 154 623 156
rect 617 152 619 154
rect 621 152 623 154
rect 617 150 623 152
rect 7 22 13 24
rect 56 22 62 24
rect 7 20 9 22
rect 11 20 13 22
rect 7 18 13 20
rect 56 20 58 22
rect 60 20 62 22
rect 56 18 62 20
rect 96 22 102 24
rect 96 20 98 22
rect 100 20 102 22
rect 96 18 102 20
rect 170 22 176 24
rect 170 20 172 22
rect 174 20 176 22
rect 170 18 176 20
rect 210 22 216 24
rect 210 20 212 22
rect 214 20 216 22
rect 210 18 216 20
rect 309 22 315 24
rect 309 20 311 22
rect 313 20 315 22
rect 309 18 315 20
rect 523 22 529 24
rect 523 20 525 22
rect 527 20 529 22
rect 523 18 529 20
rect 617 22 623 24
rect 617 20 619 22
rect 621 20 623 22
rect 617 18 623 20
<< ntie >>
rect 7 94 13 96
rect 7 92 9 94
rect 11 92 13 94
rect 56 94 62 96
rect 7 90 13 92
rect 56 92 58 94
rect 60 92 62 94
rect 129 94 135 96
rect 56 90 62 92
rect 129 92 131 94
rect 133 92 135 94
rect 170 94 176 96
rect 129 90 135 92
rect 170 92 172 94
rect 174 92 176 94
rect 243 94 249 96
rect 170 90 176 92
rect 243 92 245 94
rect 247 92 249 94
rect 309 94 315 96
rect 243 90 249 92
rect 309 92 311 94
rect 313 92 315 94
rect 523 94 529 96
rect 309 90 315 92
rect 523 92 525 94
rect 527 92 529 94
rect 584 94 590 96
rect 523 90 529 92
rect 584 92 586 94
rect 588 92 590 94
rect 584 90 590 92
rect 7 82 13 84
rect 7 80 9 82
rect 11 80 13 82
rect 56 82 62 84
rect 7 78 13 80
rect 56 80 58 82
rect 60 80 62 82
rect 129 82 135 84
rect 56 78 62 80
rect 129 80 131 82
rect 133 80 135 82
rect 170 82 176 84
rect 129 78 135 80
rect 170 80 172 82
rect 174 80 176 82
rect 243 82 249 84
rect 170 78 176 80
rect 243 80 245 82
rect 247 80 249 82
rect 309 82 315 84
rect 243 78 249 80
rect 309 80 311 82
rect 313 80 315 82
rect 523 82 529 84
rect 309 78 315 80
rect 523 80 525 82
rect 527 80 529 82
rect 584 82 590 84
rect 523 78 529 80
rect 584 80 586 82
rect 588 80 590 82
rect 584 78 590 80
<< nmos >>
rect 13 133 15 142
rect 23 133 25 139
rect 33 133 35 139
rect 62 135 64 144
rect 75 135 77 146
rect 82 135 84 146
rect 102 133 104 142
rect 118 138 120 147
rect 128 138 130 147
rect 138 138 140 150
rect 145 138 147 150
rect 176 135 178 144
rect 189 135 191 146
rect 196 135 198 146
rect 216 133 218 142
rect 232 138 234 147
rect 242 138 244 147
rect 252 138 254 150
rect 259 138 261 150
rect 287 135 289 146
rect 294 135 296 146
rect 307 135 309 144
rect 329 139 331 145
rect 339 139 341 147
rect 346 139 348 147
rect 356 139 358 147
rect 363 139 365 147
rect 373 138 375 147
rect 396 138 398 147
rect 406 139 408 147
rect 413 139 415 147
rect 423 139 425 147
rect 430 139 432 147
rect 440 139 442 145
rect 463 138 465 147
rect 473 139 475 147
rect 480 139 482 147
rect 490 139 492 147
rect 497 139 499 147
rect 507 139 509 145
rect 529 133 531 142
rect 539 133 541 139
rect 549 133 551 139
rect 572 138 574 150
rect 579 138 581 150
rect 589 138 591 147
rect 599 138 601 147
rect 615 133 617 142
rect 13 32 15 41
rect 23 35 25 41
rect 33 35 35 41
rect 62 30 64 39
rect 75 28 77 39
rect 82 28 84 39
rect 102 32 104 41
rect 118 27 120 36
rect 128 27 130 36
rect 138 24 140 36
rect 145 24 147 36
rect 176 30 178 39
rect 189 28 191 39
rect 196 28 198 39
rect 216 32 218 41
rect 232 27 234 36
rect 242 27 244 36
rect 252 24 254 36
rect 259 24 261 36
rect 287 28 289 39
rect 294 28 296 39
rect 307 30 309 39
rect 329 29 331 35
rect 339 27 341 35
rect 346 27 348 35
rect 356 27 358 35
rect 363 27 365 35
rect 373 27 375 36
rect 396 27 398 36
rect 406 27 408 35
rect 413 27 415 35
rect 423 27 425 35
rect 430 27 432 35
rect 440 29 442 35
rect 463 27 465 36
rect 473 27 475 35
rect 480 27 482 35
rect 490 27 492 35
rect 497 27 499 35
rect 507 29 509 35
rect 529 32 531 41
rect 539 35 541 41
rect 549 35 551 41
rect 572 24 574 36
rect 579 24 581 36
rect 589 27 591 36
rect 599 27 601 36
rect 615 32 617 41
<< pmos >>
rect 13 103 15 121
rect 26 93 28 114
rect 33 93 35 114
rect 62 102 64 120
rect 72 100 74 113
rect 82 100 84 113
rect 110 93 112 120
rect 126 102 128 120
rect 136 102 138 120
rect 146 93 148 120
rect 176 102 178 120
rect 186 100 188 113
rect 196 100 198 113
rect 224 93 226 120
rect 240 102 242 120
rect 250 102 252 120
rect 260 93 262 120
rect 287 100 289 113
rect 297 100 299 113
rect 307 102 309 120
rect 329 113 331 121
rect 339 93 341 109
rect 346 93 348 109
rect 356 93 358 109
rect 363 93 365 109
rect 373 93 375 111
rect 396 93 398 111
rect 440 113 442 121
rect 406 93 408 109
rect 413 93 415 109
rect 423 93 425 109
rect 430 93 432 109
rect 463 93 465 111
rect 507 113 509 121
rect 473 93 475 109
rect 480 93 482 109
rect 490 93 492 109
rect 497 93 499 109
rect 529 103 531 121
rect 542 93 544 114
rect 549 93 551 114
rect 571 93 573 120
rect 581 102 583 120
rect 591 102 593 120
rect 607 93 609 120
rect 13 53 15 71
rect 26 60 28 81
rect 33 60 35 81
rect 62 54 64 72
rect 72 61 74 74
rect 82 61 84 74
rect 110 54 112 81
rect 126 54 128 72
rect 136 54 138 72
rect 146 54 148 81
rect 176 54 178 72
rect 186 61 188 74
rect 196 61 198 74
rect 224 54 226 81
rect 240 54 242 72
rect 250 54 252 72
rect 260 54 262 81
rect 287 61 289 74
rect 297 61 299 74
rect 307 54 309 72
rect 339 65 341 81
rect 346 65 348 81
rect 356 65 358 81
rect 363 65 365 81
rect 329 53 331 61
rect 373 63 375 81
rect 396 63 398 81
rect 406 65 408 81
rect 413 65 415 81
rect 423 65 425 81
rect 430 65 432 81
rect 463 63 465 81
rect 473 65 475 81
rect 480 65 482 81
rect 490 65 492 81
rect 497 65 499 81
rect 440 53 442 61
rect 507 53 509 61
rect 529 53 531 71
rect 542 60 544 81
rect 549 60 551 81
rect 571 54 573 81
rect 581 54 583 72
rect 591 54 593 72
rect 607 54 609 81
<< polyct0 >>
rect 15 126 17 128
rect 64 126 66 128
rect 134 126 136 128
rect 144 125 146 127
rect 178 126 180 128
rect 248 126 250 128
rect 258 125 260 127
rect 305 126 307 128
rect 354 132 356 134
rect 372 131 374 133
rect 397 131 399 133
rect 347 116 349 118
rect 415 132 417 134
rect 422 116 424 118
rect 464 131 466 133
rect 482 132 484 134
rect 489 116 491 118
rect 531 126 533 128
rect 573 125 575 127
rect 583 126 585 128
rect 15 46 17 48
rect 64 46 66 48
rect 134 46 136 48
rect 144 47 146 49
rect 178 46 180 48
rect 248 46 250 48
rect 258 47 260 49
rect 305 46 307 48
rect 347 56 349 58
rect 354 40 356 42
rect 422 56 424 58
rect 372 41 374 43
rect 397 41 399 43
rect 415 40 417 42
rect 489 56 491 58
rect 464 41 466 43
rect 482 40 484 42
rect 531 46 533 48
rect 573 47 575 49
rect 583 46 585 48
<< polyct1 >>
rect 25 126 27 128
rect 74 126 76 128
rect 35 119 37 121
rect 113 131 115 133
rect 84 118 86 120
rect 188 126 190 128
rect 97 118 99 120
rect 227 131 229 133
rect 198 118 200 120
rect 295 126 297 128
rect 211 118 213 120
rect 285 118 287 120
rect 337 126 339 128
rect 364 121 366 123
rect 405 121 407 123
rect 432 126 434 128
rect 324 106 326 108
rect 472 121 474 123
rect 499 126 501 128
rect 445 106 447 108
rect 541 126 543 128
rect 512 106 514 108
rect 604 131 606 133
rect 551 119 553 121
rect 620 118 622 120
rect 35 53 37 55
rect 25 46 27 48
rect 84 54 86 56
rect 97 54 99 56
rect 74 46 76 48
rect 198 54 200 56
rect 211 54 213 56
rect 285 54 287 56
rect 113 41 115 43
rect 188 46 190 48
rect 227 41 229 43
rect 324 66 326 68
rect 295 46 297 48
rect 445 66 447 68
rect 337 46 339 48
rect 364 51 366 53
rect 405 51 407 53
rect 512 66 514 68
rect 432 46 434 48
rect 472 51 474 53
rect 499 46 501 48
rect 551 53 553 55
rect 620 54 622 56
rect 541 46 543 48
rect 604 41 606 43
<< ndifct0 >>
rect 19 148 21 150
rect 38 148 40 150
rect 28 135 30 137
rect 87 142 89 144
rect 111 143 113 145
rect 97 135 99 137
rect 123 140 125 142
rect 201 142 203 144
rect 225 143 227 145
rect 211 135 213 137
rect 237 140 239 142
rect 282 142 284 144
rect 324 141 326 143
rect 334 141 336 143
rect 351 143 353 145
rect 368 143 370 145
rect 401 143 403 145
rect 418 143 420 145
rect 435 141 437 143
rect 445 141 447 143
rect 468 143 470 145
rect 485 143 487 145
rect 535 148 537 150
rect 502 141 504 143
rect 512 141 514 143
rect 554 148 556 150
rect 544 135 546 137
rect 594 140 596 142
rect 606 143 608 145
rect 620 135 622 137
rect 28 37 30 39
rect 19 24 21 26
rect 97 37 99 39
rect 87 30 89 32
rect 111 29 113 31
rect 38 24 40 26
rect 123 32 125 34
rect 211 37 213 39
rect 201 30 203 32
rect 225 29 227 31
rect 237 32 239 34
rect 282 30 284 32
rect 324 31 326 33
rect 334 31 336 33
rect 351 29 353 31
rect 368 29 370 31
rect 401 29 403 31
rect 418 29 420 31
rect 435 31 437 33
rect 445 31 447 33
rect 468 29 470 31
rect 485 29 487 31
rect 502 31 504 33
rect 512 31 514 33
rect 544 37 546 39
rect 535 24 537 26
rect 554 24 556 26
rect 594 32 596 34
rect 620 37 622 39
rect 606 29 608 31
<< ndifct1 >>
rect 68 152 70 154
rect 8 135 10 137
rect 151 152 153 154
rect 182 152 184 154
rect 57 140 59 142
rect 133 142 135 144
rect 265 152 267 154
rect 301 152 303 154
rect 171 140 173 142
rect 247 142 249 144
rect 312 140 314 142
rect 378 140 380 142
rect 391 140 393 142
rect 458 140 460 142
rect 566 152 568 154
rect 524 135 526 137
rect 584 142 586 144
rect 8 37 10 39
rect 57 32 59 34
rect 133 30 135 32
rect 68 20 70 22
rect 171 32 173 34
rect 151 20 153 22
rect 247 30 249 32
rect 182 20 184 22
rect 312 32 314 34
rect 265 20 267 22
rect 301 20 303 22
rect 378 32 380 34
rect 391 32 393 34
rect 458 32 460 34
rect 524 37 526 39
rect 584 30 586 32
rect 566 20 568 22
<< ntiect1 >>
rect 9 92 11 94
rect 58 92 60 94
rect 131 92 133 94
rect 172 92 174 94
rect 245 92 247 94
rect 311 92 313 94
rect 525 92 527 94
rect 586 92 588 94
rect 9 80 11 82
rect 58 80 60 82
rect 131 80 133 82
rect 172 80 174 82
rect 245 80 247 82
rect 311 80 313 82
rect 525 80 527 82
rect 586 80 588 82
<< ptiect1 >>
rect 9 152 11 154
rect 58 152 60 154
rect 98 152 100 154
rect 172 152 174 154
rect 212 152 214 154
rect 311 152 313 154
rect 525 152 527 154
rect 619 152 621 154
rect 9 20 11 22
rect 58 20 60 22
rect 98 20 100 22
rect 172 20 174 22
rect 212 20 214 22
rect 311 20 313 22
rect 525 20 527 22
rect 619 20 621 22
<< pdifct0 >>
rect 19 95 21 97
rect 38 102 40 104
rect 105 116 107 118
rect 67 104 69 106
rect 77 109 79 111
rect 77 102 79 104
rect 87 102 89 104
rect 115 102 117 104
rect 131 116 133 118
rect 131 109 133 111
rect 115 95 117 97
rect 151 101 153 103
rect 219 116 221 118
rect 181 104 183 106
rect 191 109 193 111
rect 191 102 193 104
rect 201 102 203 104
rect 229 102 231 104
rect 245 116 247 118
rect 245 109 247 111
rect 229 95 231 97
rect 265 101 267 103
rect 282 102 284 104
rect 292 109 294 111
rect 292 102 294 104
rect 302 104 304 106
rect 324 117 326 119
rect 334 95 336 97
rect 351 105 353 107
rect 368 95 370 97
rect 445 117 447 119
rect 401 95 403 97
rect 418 105 420 107
rect 435 95 437 97
rect 512 117 514 119
rect 468 95 470 97
rect 485 105 487 107
rect 502 95 504 97
rect 535 95 537 97
rect 554 102 556 104
rect 566 101 568 103
rect 586 116 588 118
rect 586 109 588 111
rect 602 102 604 104
rect 602 95 604 97
rect 612 116 614 118
rect 19 77 21 79
rect 38 70 40 72
rect 67 68 69 70
rect 77 70 79 72
rect 77 63 79 65
rect 87 70 89 72
rect 105 56 107 58
rect 115 77 117 79
rect 115 70 117 72
rect 131 63 133 65
rect 131 56 133 58
rect 151 71 153 73
rect 181 68 183 70
rect 191 70 193 72
rect 191 63 193 65
rect 201 70 203 72
rect 219 56 221 58
rect 229 77 231 79
rect 229 70 231 72
rect 245 63 247 65
rect 245 56 247 58
rect 334 77 336 79
rect 265 71 267 73
rect 282 70 284 72
rect 292 70 294 72
rect 292 63 294 65
rect 302 68 304 70
rect 351 67 353 69
rect 368 77 370 79
rect 324 55 326 57
rect 401 77 403 79
rect 418 67 420 69
rect 435 77 437 79
rect 468 77 470 79
rect 485 67 487 69
rect 502 77 504 79
rect 535 77 537 79
rect 445 55 447 57
rect 512 55 514 57
rect 554 70 556 72
rect 566 71 568 73
rect 602 77 604 79
rect 586 63 588 65
rect 586 56 588 58
rect 602 70 604 72
rect 612 56 614 58
<< pdifct1 >>
rect 8 112 10 114
rect 8 105 10 107
rect 57 116 59 118
rect 57 109 59 111
rect 141 109 143 111
rect 171 116 173 118
rect 171 109 173 111
rect 255 109 257 111
rect 312 116 314 118
rect 312 109 314 111
rect 378 102 380 104
rect 391 102 393 104
rect 458 102 460 104
rect 524 112 526 114
rect 524 105 526 107
rect 576 109 578 111
rect 8 67 10 69
rect 8 60 10 62
rect 57 63 59 65
rect 57 56 59 58
rect 141 63 143 65
rect 171 63 173 65
rect 171 56 173 58
rect 255 63 257 65
rect 312 63 314 65
rect 312 56 314 58
rect 378 70 380 72
rect 391 70 393 72
rect 458 70 460 72
rect 524 67 526 69
rect 524 60 526 62
rect 576 63 578 65
<< alu0 >>
rect 17 150 23 151
rect 17 148 19 150
rect 21 148 23 150
rect 17 147 23 148
rect 36 150 42 151
rect 36 148 38 150
rect 40 148 42 150
rect 36 147 42 148
rect 109 145 115 151
rect 71 144 91 145
rect 71 142 87 144
rect 89 142 91 144
rect 109 143 111 145
rect 113 143 115 145
rect 109 142 115 143
rect 122 142 126 144
rect 71 141 91 142
rect 14 137 32 138
rect 14 135 28 137
rect 30 135 32 137
rect 14 134 32 135
rect 14 128 18 134
rect 14 126 15 128
rect 17 126 18 128
rect 10 105 11 116
rect 14 113 18 126
rect 33 121 39 122
rect 59 138 60 140
rect 71 137 75 141
rect 122 140 123 142
rect 125 140 126 142
rect 63 133 75 137
rect 63 128 67 133
rect 63 126 64 128
rect 66 126 67 128
rect 14 109 29 113
rect 25 105 29 109
rect 63 114 67 126
rect 96 137 100 139
rect 96 135 97 137
rect 99 135 100 137
rect 96 129 100 135
rect 122 137 126 140
rect 122 133 146 137
rect 96 125 107 129
rect 63 111 80 114
rect 63 110 77 111
rect 76 109 77 110
rect 79 109 80 111
rect 65 106 71 107
rect 25 104 42 105
rect 25 102 38 104
rect 40 102 42 104
rect 25 101 42 102
rect 65 104 67 106
rect 69 104 71 106
rect 17 97 23 98
rect 17 95 19 97
rect 21 95 23 97
rect 65 95 71 104
rect 76 104 80 109
rect 103 119 107 125
rect 142 129 146 133
rect 122 128 138 129
rect 122 126 134 128
rect 136 126 138 128
rect 122 125 138 126
rect 142 127 147 129
rect 142 125 144 127
rect 146 125 147 127
rect 122 119 126 125
rect 142 123 147 125
rect 142 121 146 123
rect 103 118 126 119
rect 103 116 105 118
rect 107 116 126 118
rect 103 115 126 116
rect 76 102 77 104
rect 79 102 80 104
rect 76 100 80 102
rect 85 104 91 105
rect 85 102 87 104
rect 89 102 91 104
rect 85 95 91 102
rect 114 104 118 106
rect 114 102 115 104
rect 117 102 118 104
rect 114 97 118 102
rect 122 104 126 115
rect 130 118 146 121
rect 130 116 131 118
rect 133 117 146 118
rect 133 116 134 117
rect 130 111 134 116
rect 130 109 131 111
rect 133 109 134 111
rect 130 107 134 109
rect 223 145 229 151
rect 185 144 205 145
rect 185 142 201 144
rect 203 142 205 144
rect 223 143 225 145
rect 227 143 229 145
rect 223 142 229 143
rect 236 142 240 144
rect 185 141 205 142
rect 173 138 174 140
rect 185 137 189 141
rect 236 140 237 142
rect 239 140 240 142
rect 280 144 300 145
rect 280 142 282 144
rect 284 142 300 144
rect 280 141 300 142
rect 177 133 189 137
rect 177 128 181 133
rect 177 126 178 128
rect 180 126 181 128
rect 177 114 181 126
rect 210 137 214 139
rect 210 135 211 137
rect 213 135 214 137
rect 210 129 214 135
rect 236 137 240 140
rect 236 133 260 137
rect 210 125 221 129
rect 217 119 221 125
rect 256 129 260 133
rect 236 128 252 129
rect 236 126 248 128
rect 250 126 252 128
rect 236 125 252 126
rect 256 127 261 129
rect 256 125 258 127
rect 260 125 261 127
rect 236 119 240 125
rect 256 123 261 125
rect 256 121 260 123
rect 217 118 240 119
rect 217 116 219 118
rect 221 116 240 118
rect 217 115 240 116
rect 177 111 194 114
rect 177 110 191 111
rect 190 109 191 110
rect 193 109 194 111
rect 179 106 185 107
rect 179 104 181 106
rect 183 104 185 106
rect 122 103 155 104
rect 122 101 151 103
rect 153 101 155 103
rect 122 100 155 101
rect 114 95 115 97
rect 117 95 118 97
rect 179 95 185 104
rect 190 104 194 109
rect 190 102 191 104
rect 193 102 194 104
rect 190 100 194 102
rect 199 104 205 105
rect 199 102 201 104
rect 203 102 205 104
rect 199 100 205 102
rect 228 104 232 106
rect 228 102 229 104
rect 231 102 232 104
rect 199 95 201 100
rect 228 97 232 102
rect 236 104 240 115
rect 244 118 260 121
rect 244 116 245 118
rect 247 117 260 118
rect 296 137 300 141
rect 311 138 312 140
rect 296 133 308 137
rect 304 128 308 133
rect 304 126 305 128
rect 307 126 308 128
rect 247 116 248 117
rect 244 111 248 116
rect 244 109 245 111
rect 247 109 248 111
rect 244 107 248 109
rect 304 114 308 126
rect 291 111 308 114
rect 291 109 292 111
rect 294 110 308 111
rect 322 143 328 144
rect 322 141 324 143
rect 326 141 328 143
rect 322 140 328 141
rect 332 143 338 151
rect 332 141 334 143
rect 336 141 338 143
rect 349 145 364 146
rect 349 143 351 145
rect 353 143 364 145
rect 349 142 364 143
rect 332 140 338 141
rect 322 120 326 140
rect 360 137 364 142
rect 367 145 371 151
rect 367 143 368 145
rect 370 143 371 145
rect 367 141 371 143
rect 346 134 357 136
rect 346 132 354 134
rect 356 132 357 134
rect 360 135 374 137
rect 360 133 375 135
rect 346 130 357 132
rect 370 131 372 133
rect 374 131 375 133
rect 346 120 350 130
rect 370 129 375 131
rect 322 119 350 120
rect 322 117 324 119
rect 326 118 350 119
rect 326 117 347 118
rect 322 116 347 117
rect 349 116 350 118
rect 366 119 367 125
rect 346 114 350 116
rect 294 109 295 110
rect 280 104 286 105
rect 236 103 269 104
rect 236 101 265 103
rect 267 101 269 103
rect 236 100 269 101
rect 280 102 282 104
rect 284 102 286 104
rect 228 95 229 97
rect 231 95 232 97
rect 280 95 286 102
rect 291 104 295 109
rect 370 112 374 129
rect 358 108 374 112
rect 291 102 292 104
rect 294 102 295 104
rect 291 100 295 102
rect 300 106 306 107
rect 300 104 302 106
rect 304 104 306 106
rect 300 95 306 104
rect 349 107 362 108
rect 349 105 351 107
rect 353 105 362 107
rect 349 104 362 105
rect 400 145 404 151
rect 400 143 401 145
rect 403 143 404 145
rect 400 141 404 143
rect 407 145 422 146
rect 407 143 418 145
rect 420 143 422 145
rect 407 142 422 143
rect 433 143 439 151
rect 467 145 471 151
rect 407 137 411 142
rect 433 141 435 143
rect 437 141 439 143
rect 433 140 439 141
rect 443 143 449 144
rect 443 141 445 143
rect 447 141 449 143
rect 443 140 449 141
rect 397 135 411 137
rect 396 133 411 135
rect 414 134 425 136
rect 396 131 397 133
rect 399 131 401 133
rect 396 129 401 131
rect 414 132 415 134
rect 417 132 425 134
rect 414 130 425 132
rect 397 112 401 129
rect 404 119 405 125
rect 421 120 425 130
rect 445 120 449 140
rect 421 119 449 120
rect 421 118 445 119
rect 421 116 422 118
rect 424 117 445 118
rect 447 117 449 119
rect 424 116 449 117
rect 467 143 468 145
rect 470 143 471 145
rect 467 141 471 143
rect 474 145 489 146
rect 474 143 485 145
rect 487 143 489 145
rect 474 142 489 143
rect 500 143 506 151
rect 533 150 539 151
rect 533 148 535 150
rect 537 148 539 150
rect 533 147 539 148
rect 552 150 558 151
rect 552 148 554 150
rect 556 148 558 150
rect 552 147 558 148
rect 604 145 610 151
rect 474 137 478 142
rect 500 141 502 143
rect 504 141 506 143
rect 500 140 506 141
rect 510 143 516 144
rect 510 141 512 143
rect 514 141 516 143
rect 510 140 516 141
rect 464 135 478 137
rect 421 114 425 116
rect 397 108 413 112
rect 409 107 422 108
rect 409 105 418 107
rect 420 105 422 107
rect 409 104 422 105
rect 463 133 478 135
rect 481 134 492 136
rect 463 131 464 133
rect 466 131 468 133
rect 463 129 468 131
rect 481 132 482 134
rect 484 132 492 134
rect 481 130 492 132
rect 464 112 468 129
rect 471 119 472 125
rect 488 120 492 130
rect 512 120 516 140
rect 593 142 597 144
rect 604 143 606 145
rect 608 143 610 145
rect 604 142 610 143
rect 488 119 516 120
rect 488 118 512 119
rect 488 116 489 118
rect 491 117 512 118
rect 514 117 516 119
rect 491 116 516 117
rect 530 137 548 138
rect 530 135 544 137
rect 546 135 548 137
rect 530 134 548 135
rect 488 114 492 116
rect 530 128 534 134
rect 530 126 531 128
rect 533 126 534 128
rect 464 108 480 112
rect 476 107 489 108
rect 476 105 485 107
rect 487 105 489 107
rect 476 104 489 105
rect 526 105 527 116
rect 530 113 534 126
rect 593 140 594 142
rect 596 140 597 142
rect 593 137 597 140
rect 549 121 555 122
rect 530 109 545 113
rect 541 105 545 109
rect 573 133 597 137
rect 573 129 577 133
rect 619 137 623 139
rect 619 135 620 137
rect 622 135 623 137
rect 572 127 577 129
rect 572 125 573 127
rect 575 125 577 127
rect 581 128 597 129
rect 581 126 583 128
rect 585 126 597 128
rect 581 125 597 126
rect 572 123 577 125
rect 573 121 577 123
rect 573 118 589 121
rect 573 117 586 118
rect 585 116 586 117
rect 588 116 589 118
rect 585 111 589 116
rect 585 109 586 111
rect 588 109 589 111
rect 585 107 589 109
rect 593 119 597 125
rect 619 129 623 135
rect 612 125 623 129
rect 612 119 616 125
rect 593 118 616 119
rect 593 116 612 118
rect 614 116 616 118
rect 593 115 616 116
rect 541 104 558 105
rect 593 104 597 115
rect 541 102 554 104
rect 556 102 558 104
rect 541 101 558 102
rect 564 103 597 104
rect 564 101 566 103
rect 568 101 597 103
rect 564 100 597 101
rect 601 104 605 106
rect 601 102 602 104
rect 604 102 605 104
rect 333 97 337 99
rect 333 95 334 97
rect 336 95 337 97
rect 366 97 372 98
rect 366 95 368 97
rect 370 95 372 97
rect 399 97 405 98
rect 399 95 401 97
rect 403 95 405 97
rect 434 97 438 99
rect 434 95 435 97
rect 437 95 438 97
rect 466 97 472 98
rect 466 95 468 97
rect 470 95 472 97
rect 501 97 505 99
rect 501 95 502 97
rect 504 95 505 97
rect 533 97 539 98
rect 533 95 535 97
rect 537 95 539 97
rect 601 97 605 102
rect 601 95 602 97
rect 604 95 605 97
rect 17 77 19 79
rect 21 77 23 79
rect 17 76 23 77
rect 25 72 42 73
rect 25 70 38 72
rect 40 70 42 72
rect 25 69 42 70
rect 65 70 71 79
rect 10 58 11 69
rect 25 65 29 69
rect 65 68 67 70
rect 69 68 71 70
rect 65 67 71 68
rect 76 72 80 74
rect 76 70 77 72
rect 79 70 80 72
rect 14 61 29 65
rect 76 65 80 70
rect 85 72 91 79
rect 114 77 115 79
rect 117 77 118 79
rect 85 70 87 72
rect 89 70 91 72
rect 85 69 91 70
rect 114 72 118 77
rect 114 70 115 72
rect 117 70 118 72
rect 114 68 118 70
rect 122 73 155 74
rect 122 71 151 73
rect 153 71 155 73
rect 122 70 155 71
rect 179 70 185 79
rect 76 64 77 65
rect 14 48 18 61
rect 63 63 77 64
rect 79 63 80 65
rect 63 60 80 63
rect 33 52 39 53
rect 14 46 15 48
rect 17 46 18 48
rect 14 40 18 46
rect 14 39 32 40
rect 14 37 28 39
rect 30 37 32 39
rect 14 36 32 37
rect 63 48 67 60
rect 122 59 126 70
rect 179 68 181 70
rect 183 68 185 70
rect 179 67 185 68
rect 190 72 194 74
rect 190 70 191 72
rect 193 70 194 72
rect 103 58 126 59
rect 103 56 105 58
rect 107 56 126 58
rect 103 55 126 56
rect 103 49 107 55
rect 63 46 64 48
rect 66 46 67 48
rect 63 41 67 46
rect 63 37 75 41
rect 59 34 60 36
rect 71 33 75 37
rect 96 45 107 49
rect 96 39 100 45
rect 122 49 126 55
rect 130 65 134 67
rect 130 63 131 65
rect 133 63 134 65
rect 130 58 134 63
rect 130 56 131 58
rect 133 57 134 58
rect 133 56 146 57
rect 130 53 146 56
rect 142 51 146 53
rect 142 49 147 51
rect 122 48 138 49
rect 122 46 134 48
rect 136 46 138 48
rect 122 45 138 46
rect 142 47 144 49
rect 146 47 147 49
rect 142 45 147 47
rect 96 37 97 39
rect 99 37 100 39
rect 96 35 100 37
rect 142 41 146 45
rect 122 37 146 41
rect 122 34 126 37
rect 71 32 91 33
rect 122 32 123 34
rect 125 32 126 34
rect 71 30 87 32
rect 89 30 91 32
rect 71 29 91 30
rect 109 31 115 32
rect 109 29 111 31
rect 113 29 115 31
rect 122 30 126 32
rect 190 65 194 70
rect 199 72 205 79
rect 228 77 229 79
rect 231 77 232 79
rect 199 70 201 72
rect 203 70 205 72
rect 199 69 205 70
rect 228 72 232 77
rect 228 70 229 72
rect 231 70 232 72
rect 228 68 232 70
rect 236 73 269 74
rect 236 71 265 73
rect 267 71 269 73
rect 236 70 269 71
rect 280 72 286 79
rect 280 70 282 72
rect 284 70 286 72
rect 190 64 191 65
rect 177 63 191 64
rect 193 63 194 65
rect 177 60 194 63
rect 177 48 181 60
rect 236 59 240 70
rect 280 69 286 70
rect 291 72 295 74
rect 291 70 292 72
rect 294 70 295 72
rect 217 58 240 59
rect 217 56 219 58
rect 221 56 240 58
rect 217 55 240 56
rect 217 49 221 55
rect 177 46 178 48
rect 180 46 181 48
rect 177 41 181 46
rect 177 37 189 41
rect 173 34 174 36
rect 17 26 23 27
rect 17 24 19 26
rect 21 24 23 26
rect 17 23 23 24
rect 36 26 42 27
rect 36 24 38 26
rect 40 24 42 26
rect 36 23 42 24
rect 109 23 115 29
rect 185 33 189 37
rect 210 45 221 49
rect 210 39 214 45
rect 236 49 240 55
rect 244 65 248 67
rect 244 63 245 65
rect 247 63 248 65
rect 244 58 248 63
rect 244 56 245 58
rect 247 57 248 58
rect 247 56 260 57
rect 244 53 260 56
rect 256 51 260 53
rect 291 65 295 70
rect 300 70 306 79
rect 333 77 334 79
rect 336 77 337 79
rect 333 75 337 77
rect 366 77 368 79
rect 370 77 372 79
rect 366 76 372 77
rect 399 77 401 79
rect 403 77 405 79
rect 399 76 405 77
rect 434 77 435 79
rect 437 77 438 79
rect 434 75 438 77
rect 466 77 468 79
rect 470 77 472 79
rect 466 76 472 77
rect 501 77 502 79
rect 504 77 505 79
rect 501 75 505 77
rect 533 77 535 79
rect 537 77 539 79
rect 533 76 539 77
rect 601 77 602 79
rect 604 77 605 79
rect 300 68 302 70
rect 304 68 306 70
rect 300 67 306 68
rect 291 63 292 65
rect 294 64 295 65
rect 294 63 308 64
rect 291 60 308 63
rect 256 49 261 51
rect 236 48 252 49
rect 236 46 248 48
rect 250 46 252 48
rect 236 45 252 46
rect 256 47 258 49
rect 260 47 261 49
rect 256 45 261 47
rect 210 37 211 39
rect 213 37 214 39
rect 210 35 214 37
rect 256 41 260 45
rect 236 37 260 41
rect 236 34 240 37
rect 185 32 205 33
rect 236 32 237 34
rect 239 32 240 34
rect 304 48 308 60
rect 349 69 362 70
rect 349 67 351 69
rect 353 67 362 69
rect 349 66 362 67
rect 358 62 374 66
rect 346 58 350 60
rect 304 46 305 48
rect 307 46 308 48
rect 304 41 308 46
rect 296 37 308 41
rect 296 33 300 37
rect 311 34 312 36
rect 185 30 201 32
rect 203 30 205 32
rect 185 29 205 30
rect 223 31 229 32
rect 223 29 225 31
rect 227 29 229 31
rect 236 30 240 32
rect 280 32 300 33
rect 280 30 282 32
rect 284 30 300 32
rect 280 29 300 30
rect 223 23 229 29
rect 322 57 347 58
rect 322 55 324 57
rect 326 56 347 57
rect 349 56 350 58
rect 326 55 350 56
rect 322 54 350 55
rect 322 34 326 54
rect 346 44 350 54
rect 366 49 367 55
rect 370 45 374 62
rect 346 42 357 44
rect 346 40 354 42
rect 356 40 357 42
rect 370 43 375 45
rect 370 41 372 43
rect 374 41 375 43
rect 346 38 357 40
rect 360 39 375 41
rect 360 37 374 39
rect 322 33 328 34
rect 322 31 324 33
rect 326 31 328 33
rect 322 30 328 31
rect 332 33 338 34
rect 332 31 334 33
rect 336 31 338 33
rect 360 32 364 37
rect 332 23 338 31
rect 349 31 364 32
rect 349 29 351 31
rect 353 29 364 31
rect 349 28 364 29
rect 367 31 371 33
rect 367 29 368 31
rect 370 29 371 31
rect 367 23 371 29
rect 409 69 422 70
rect 409 67 418 69
rect 420 67 422 69
rect 409 66 422 67
rect 397 62 413 66
rect 397 45 401 62
rect 476 69 489 70
rect 421 58 425 60
rect 404 49 405 55
rect 421 56 422 58
rect 424 57 449 58
rect 424 56 445 57
rect 421 55 445 56
rect 447 55 449 57
rect 421 54 449 55
rect 396 43 401 45
rect 421 44 425 54
rect 396 41 397 43
rect 399 41 401 43
rect 414 42 425 44
rect 396 39 411 41
rect 397 37 411 39
rect 414 40 415 42
rect 417 40 425 42
rect 414 38 425 40
rect 400 31 404 33
rect 400 29 401 31
rect 403 29 404 31
rect 400 23 404 29
rect 407 32 411 37
rect 445 34 449 54
rect 433 33 439 34
rect 407 31 422 32
rect 407 29 418 31
rect 420 29 422 31
rect 407 28 422 29
rect 433 31 435 33
rect 437 31 439 33
rect 433 23 439 31
rect 443 33 449 34
rect 443 31 445 33
rect 447 31 449 33
rect 443 30 449 31
rect 476 67 485 69
rect 487 67 489 69
rect 476 66 489 67
rect 464 62 480 66
rect 464 45 468 62
rect 564 73 597 74
rect 541 72 558 73
rect 541 70 554 72
rect 556 70 558 72
rect 564 71 566 73
rect 568 71 597 73
rect 564 70 597 71
rect 541 69 558 70
rect 488 58 492 60
rect 471 49 472 55
rect 488 56 489 58
rect 491 57 516 58
rect 491 56 512 57
rect 488 55 512 56
rect 514 55 516 57
rect 488 54 516 55
rect 463 43 468 45
rect 488 44 492 54
rect 463 41 464 43
rect 466 41 468 43
rect 481 42 492 44
rect 463 39 478 41
rect 464 37 478 39
rect 481 40 482 42
rect 484 40 492 42
rect 481 38 492 40
rect 467 31 471 33
rect 467 29 468 31
rect 470 29 471 31
rect 467 23 471 29
rect 474 32 478 37
rect 512 34 516 54
rect 526 58 527 69
rect 541 65 545 69
rect 530 61 545 65
rect 530 48 534 61
rect 585 65 589 67
rect 585 63 586 65
rect 588 63 589 65
rect 549 52 555 53
rect 530 46 531 48
rect 533 46 534 48
rect 530 40 534 46
rect 530 39 548 40
rect 530 37 544 39
rect 546 37 548 39
rect 530 36 548 37
rect 585 58 589 63
rect 585 57 586 58
rect 573 56 586 57
rect 588 56 589 58
rect 573 53 589 56
rect 593 59 597 70
rect 601 72 605 77
rect 601 70 602 72
rect 604 70 605 72
rect 601 68 605 70
rect 593 58 616 59
rect 593 56 612 58
rect 614 56 616 58
rect 593 55 616 56
rect 573 51 577 53
rect 572 49 577 51
rect 593 49 597 55
rect 572 47 573 49
rect 575 47 577 49
rect 572 45 577 47
rect 581 48 597 49
rect 581 46 583 48
rect 585 46 597 48
rect 581 45 597 46
rect 500 33 506 34
rect 474 31 489 32
rect 474 29 485 31
rect 487 29 489 31
rect 474 28 489 29
rect 500 31 502 33
rect 504 31 506 33
rect 500 23 506 31
rect 510 33 516 34
rect 510 31 512 33
rect 514 31 516 33
rect 510 30 516 31
rect 573 41 577 45
rect 612 49 616 55
rect 612 45 623 49
rect 573 37 597 41
rect 593 34 597 37
rect 619 39 623 45
rect 619 37 620 39
rect 622 37 623 39
rect 619 35 623 37
rect 593 32 594 34
rect 596 32 597 34
rect 593 30 597 32
rect 604 31 610 32
rect 604 29 606 31
rect 608 29 610 31
rect 533 26 539 27
rect 533 24 535 26
rect 537 24 539 26
rect 533 23 539 24
rect 552 26 558 27
rect 552 24 554 26
rect 556 24 558 26
rect 552 23 558 24
rect 604 23 610 29
<< via1 >>
rect 39 126 41 128
rect 80 135 82 137
rect 105 135 107 137
rect 88 111 90 113
rect 152 134 154 136
rect 97 111 99 113
rect 170 126 172 128
rect 194 135 196 137
rect 219 135 221 137
rect 202 111 204 113
rect 211 111 213 113
rect 211 102 213 104
rect 266 119 268 121
rect 313 134 315 136
rect 330 134 332 136
rect 355 118 357 120
rect 332 110 334 112
rect 379 126 381 128
rect 406 126 408 128
rect 437 134 439 136
rect 457 134 459 136
rect 480 119 482 121
rect 505 134 507 136
rect 523 118 525 120
rect 504 110 506 112
rect 565 134 567 136
rect 7 55 9 57
rect 88 61 90 63
rect 39 46 41 48
rect 97 61 99 63
rect 80 37 82 39
rect 105 37 107 39
rect 152 38 154 40
rect 202 61 204 63
rect 170 46 172 48
rect 211 61 213 63
rect 194 37 196 39
rect 266 53 268 55
rect 219 37 221 39
rect 332 62 334 64
rect 313 38 315 40
rect 330 38 332 40
rect 355 54 357 56
rect 379 46 381 48
rect 406 46 408 48
rect 437 38 439 40
rect 504 62 506 64
rect 480 53 482 55
rect 457 38 459 40
rect 505 38 507 40
rect 523 54 525 56
rect 565 38 567 40
<< labels >>
rlabel alu1 125 155 125 155 8 vss
rlabel alu1 125 91 125 91 8 vdd
rlabel alu1 73 91 73 91 8 vdd
rlabel alu1 73 155 73 155 8 vss
rlabel alu1 239 155 239 155 8 vss
rlabel alu1 239 91 239 91 8 vdd
rlabel alu1 187 91 187 91 8 vdd
rlabel alu1 187 155 187 155 8 vss
rlabel alu1 24 155 24 155 8 vss
rlabel alu1 24 91 24 91 8 vdd
rlabel alu1 298 155 298 155 2 vss
rlabel alu1 298 91 298 91 2 vdd
rlabel alu1 419 155 419 155 8 vss
rlabel alu1 419 91 419 91 8 vdd
rlabel alu1 352 155 352 155 2 vss
rlabel alu1 352 91 352 91 2 vdd
rlabel alu1 486 155 486 155 8 vss
rlabel alu1 486 91 486 91 8 vdd
rlabel alu1 540 155 540 155 8 vss
rlabel alu1 540 91 540 91 8 vdd
rlabel alu1 594 155 594 155 2 vss
rlabel alu1 594 91 594 91 2 vdd
rlabel alu1 8 125 8 125 1 cout2
rlabel alu2 73 128 73 128 1 a1
rlabel via1 88 113 88 113 1 b1
rlabel alu1 290 131 290 131 1 a1
rlabel alu1 298 127 298 127 1 a1
rlabel alu1 282 111 282 111 1 b1
rlabel alu1 399 103 399 103 1 z1
rlabel alu1 540 127 540 127 1 a1
rlabel alu1 548 127 548 127 1 a1
rlabel alu1 540 119 540 119 1 b1
rlabel alu1 548 119 548 119 1 b1
rlabel alu1 556 111 556 111 1 b1
rlabel alu1 614 103 614 103 1 b1
rlabel alu1 622 111 622 111 1 b1
rlabel polyct1 606 131 606 131 1 a1
rlabel alu1 614 135 614 135 1 a1
rlabel alu1 391 122 391 122 1 z1
rlabel alu1 125 19 125 19 6 vss
rlabel alu1 125 83 125 83 6 vdd
rlabel alu1 73 83 73 83 6 vdd
rlabel alu1 73 19 73 19 6 vss
rlabel alu1 239 19 239 19 6 vss
rlabel alu1 239 83 239 83 6 vdd
rlabel alu1 187 83 187 83 6 vdd
rlabel alu1 187 19 187 19 6 vss
rlabel alu1 24 19 24 19 6 vss
rlabel alu1 24 83 24 83 6 vdd
rlabel via1 204 62 204 62 1 cin
rlabel alu1 298 19 298 19 4 vss
rlabel alu1 298 83 298 83 4 vdd
rlabel alu1 419 19 419 19 6 vss
rlabel alu1 419 83 419 83 6 vdd
rlabel alu1 352 19 352 19 4 vss
rlabel alu1 352 83 352 83 4 vdd
rlabel alu1 486 19 486 19 6 vss
rlabel alu1 486 83 486 83 6 vdd
rlabel alu1 540 19 540 19 6 vss
rlabel alu1 540 83 540 83 6 vdd
rlabel alu1 594 19 594 19 4 vss
rlabel alu1 594 83 594 83 4 vdd
rlabel alu2 73 46 73 46 1 a0
rlabel via1 88 61 88 61 1 b0
rlabel alu1 290 43 290 43 1 a0
rlabel alu1 298 47 298 47 1 a0
rlabel alu1 282 63 282 63 1 b0
rlabel alu1 391 52 391 52 1 z0
rlabel alu1 548 47 548 47 1 a0
rlabel alu1 540 47 540 47 1 a0
rlabel alu1 540 55 540 55 1 b0
rlabel alu1 548 55 548 55 1 b0
rlabel alu1 556 63 556 63 1 b0
rlabel polyct1 606 43 606 43 1 a0
rlabel alu1 614 39 614 39 1 a0
rlabel alu1 614 71 614 71 1 b0
rlabel alu1 622 63 622 63 1 b0
rlabel alu1 399 71 399 71 1 z0
rlabel alu1 8 48 8 48 1 cout1
rlabel alu1 447 71 447 71 1 s00
rlabel alu1 324 71 324 71 1 s01
rlabel via1 332 63 332 63 1 s01
rlabel alu1 514 71 514 71 1 s01
rlabel via1 506 63 506 63 1 s01
rlabel alu1 447 103 447 103 1 s10
rlabel alu1 514 103 514 103 1 s11
rlabel via1 506 111 506 111 1 s11
rlabel alu1 324 103 324 103 1 s11
rlabel via1 332 111 332 111 1 s11
rlabel via1 212 103 212 103 1 cout1
rlabel via1 203 112 203 112 1 cout1
<< end >>
