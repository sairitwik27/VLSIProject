magic
tech scmos
timestamp 1607761418
<< ab >>
rect 88 323 94 328
rect 202 323 208 328
rect 4 35 44 323
rect 53 291 157 323
rect 53 259 93 291
rect 94 259 157 291
rect 46 243 51 259
rect 53 243 157 259
rect 53 211 93 243
rect 94 211 157 243
rect 53 147 157 211
rect 53 115 93 147
rect 94 115 157 147
rect 46 99 51 115
rect 53 99 157 115
rect 53 67 93 99
rect 94 67 157 99
rect 53 35 157 67
rect 167 291 271 323
rect 272 315 276 323
rect 167 259 207 291
rect 208 259 271 291
rect 167 243 271 259
rect 272 243 274 259
rect 167 211 207 243
rect 208 211 271 243
rect 167 147 271 211
rect 272 171 276 187
rect 167 115 207 147
rect 208 115 271 147
rect 167 99 271 115
rect 272 99 274 115
rect 167 67 207 99
rect 208 67 271 99
rect 167 35 271 67
rect 272 35 276 43
rect 278 35 318 323
rect 319 315 383 323
rect 322 259 383 315
rect 319 243 383 259
rect 322 187 383 243
rect 319 171 383 187
rect 322 115 383 171
rect 319 99 383 115
rect 322 43 383 99
rect 319 35 383 43
rect 387 35 451 323
rect 455 35 518 323
rect 520 315 560 323
rect 562 315 632 323
rect 521 259 560 315
rect 563 259 626 315
rect 520 243 560 259
rect 561 243 626 259
rect 627 243 632 259
rect 521 187 560 243
rect 563 187 626 243
rect 520 171 560 187
rect 562 171 632 187
rect 521 115 560 171
rect 563 115 626 171
rect 520 99 560 115
rect 561 99 626 115
rect 627 99 632 115
rect 521 43 560 99
rect 563 43 626 99
rect 520 35 560 43
rect 562 35 632 43
rect 88 30 94 35
rect 202 30 208 35
<< nwell >>
rect -1 211 632 291
rect -1 67 632 147
<< pwell >>
rect -1 291 632 328
rect -1 147 632 211
rect -1 30 632 67
<< poly >>
rect 13 306 15 311
rect 23 303 25 308
rect 33 303 35 308
rect 62 308 64 312
rect 75 310 77 315
rect 82 310 84 315
rect 105 319 130 321
rect 105 311 107 319
rect 118 311 120 315
rect 128 311 130 319
rect 138 314 140 319
rect 145 314 147 319
rect 102 309 107 311
rect 102 306 104 309
rect 13 294 15 297
rect 23 294 25 297
rect 13 292 19 294
rect 13 290 15 292
rect 17 290 19 292
rect 13 288 19 290
rect 23 292 29 294
rect 23 290 25 292
rect 27 290 29 292
rect 23 288 29 290
rect 13 285 15 288
rect 26 278 28 288
rect 33 287 35 297
rect 62 294 64 299
rect 75 294 77 299
rect 62 292 68 294
rect 62 290 64 292
rect 66 290 68 292
rect 62 288 68 290
rect 72 292 78 294
rect 72 290 74 292
rect 76 290 78 292
rect 72 288 78 290
rect 33 285 39 287
rect 33 283 35 285
rect 37 283 39 285
rect 62 284 64 288
rect 33 281 39 283
rect 33 278 35 281
rect 13 262 15 267
rect 72 277 74 288
rect 82 286 84 299
rect 176 308 178 312
rect 189 310 191 315
rect 196 310 198 315
rect 219 319 244 321
rect 219 311 221 319
rect 232 311 234 315
rect 242 311 244 319
rect 252 314 254 319
rect 259 314 261 319
rect 118 299 120 302
rect 111 297 120 299
rect 128 298 130 302
rect 138 299 140 302
rect 102 289 104 297
rect 111 295 113 297
rect 115 295 120 297
rect 111 293 120 295
rect 136 297 140 299
rect 136 294 138 297
rect 118 289 120 293
rect 132 292 138 294
rect 145 293 147 302
rect 216 309 221 311
rect 216 306 218 309
rect 176 294 178 299
rect 189 294 191 299
rect 132 290 134 292
rect 136 290 138 292
rect 99 287 112 289
rect 118 287 128 289
rect 132 288 138 290
rect 99 286 101 287
rect 82 284 88 286
rect 82 282 84 284
rect 86 282 88 284
rect 82 280 88 282
rect 95 284 101 286
rect 110 284 112 287
rect 126 284 128 287
rect 136 284 138 288
rect 142 291 148 293
rect 142 289 144 291
rect 146 289 148 291
rect 142 287 148 289
rect 146 284 148 287
rect 176 292 182 294
rect 176 290 178 292
rect 180 290 182 292
rect 176 288 182 290
rect 186 292 192 294
rect 186 290 188 292
rect 190 290 192 292
rect 186 288 192 290
rect 176 284 178 288
rect 95 282 97 284
rect 99 282 101 284
rect 95 280 101 282
rect 82 277 84 280
rect 62 262 64 266
rect 72 259 74 264
rect 82 259 84 264
rect 26 253 28 257
rect 33 253 35 257
rect 126 262 128 266
rect 136 262 138 266
rect 110 253 112 257
rect 186 277 188 288
rect 196 286 198 299
rect 287 310 289 315
rect 294 310 296 315
rect 329 319 348 321
rect 232 299 234 302
rect 225 297 234 299
rect 242 298 244 302
rect 252 299 254 302
rect 216 289 218 297
rect 225 295 227 297
rect 229 295 234 297
rect 225 293 234 295
rect 250 297 254 299
rect 250 294 252 297
rect 232 289 234 293
rect 246 292 252 294
rect 259 293 261 302
rect 307 308 309 312
rect 329 309 331 319
rect 339 311 341 315
rect 346 311 348 319
rect 423 319 442 321
rect 356 311 358 316
rect 363 311 365 316
rect 373 311 375 316
rect 396 311 398 316
rect 406 311 408 316
rect 413 311 415 316
rect 423 311 425 319
rect 430 311 432 315
rect 246 290 248 292
rect 250 290 252 292
rect 213 287 226 289
rect 232 287 242 289
rect 246 288 252 290
rect 213 286 215 287
rect 196 284 202 286
rect 196 282 198 284
rect 200 282 202 284
rect 196 280 202 282
rect 209 284 215 286
rect 224 284 226 287
rect 240 284 242 287
rect 250 284 252 288
rect 256 291 262 293
rect 256 289 258 291
rect 260 289 262 291
rect 256 287 262 289
rect 260 284 262 287
rect 287 286 289 299
rect 294 294 296 299
rect 307 294 309 299
rect 293 292 299 294
rect 293 290 295 292
rect 297 290 299 292
rect 293 288 299 290
rect 303 292 309 294
rect 303 290 305 292
rect 307 290 309 292
rect 303 288 309 290
rect 283 284 289 286
rect 209 282 211 284
rect 213 282 215 284
rect 209 280 215 282
rect 196 277 198 280
rect 176 262 178 266
rect 186 259 188 264
rect 196 259 198 264
rect 146 253 148 257
rect 240 262 242 266
rect 250 262 252 266
rect 224 253 226 257
rect 283 282 285 284
rect 287 282 289 284
rect 283 280 289 282
rect 287 277 289 280
rect 297 277 299 288
rect 307 284 309 288
rect 329 285 331 303
rect 339 294 341 303
rect 335 292 341 294
rect 335 290 337 292
rect 339 290 341 292
rect 335 288 341 290
rect 346 290 348 303
rect 356 300 358 303
rect 352 298 358 300
rect 352 296 354 298
rect 356 296 358 298
rect 352 294 358 296
rect 346 288 358 290
rect 363 289 365 303
rect 440 309 442 319
rect 490 319 509 321
rect 463 311 465 316
rect 473 311 475 316
rect 480 311 482 316
rect 490 311 492 319
rect 497 311 499 315
rect 373 299 375 302
rect 396 299 398 302
rect 370 297 376 299
rect 370 295 372 297
rect 374 295 376 297
rect 370 293 376 295
rect 395 297 401 299
rect 395 295 397 297
rect 399 295 401 297
rect 395 293 401 295
rect 329 274 331 277
rect 322 272 331 274
rect 339 273 341 288
rect 345 282 351 284
rect 345 280 347 282
rect 349 280 351 282
rect 345 278 351 280
rect 346 273 348 278
rect 356 273 358 288
rect 362 287 368 289
rect 362 285 364 287
rect 366 285 368 287
rect 362 283 368 285
rect 363 273 365 283
rect 373 275 375 293
rect 396 275 398 293
rect 406 289 408 303
rect 413 300 415 303
rect 413 298 419 300
rect 413 296 415 298
rect 417 296 419 298
rect 413 294 419 296
rect 423 290 425 303
rect 403 287 409 289
rect 403 285 405 287
rect 407 285 409 287
rect 403 283 409 285
rect 413 288 425 290
rect 430 294 432 303
rect 430 292 436 294
rect 430 290 432 292
rect 434 290 436 292
rect 430 288 436 290
rect 322 270 324 272
rect 326 270 328 272
rect 322 268 328 270
rect 287 259 289 264
rect 297 259 299 264
rect 307 262 309 266
rect 260 253 262 257
rect 406 273 408 283
rect 413 273 415 288
rect 420 282 426 284
rect 420 280 422 282
rect 424 280 426 282
rect 420 278 426 280
rect 423 273 425 278
rect 430 273 432 288
rect 440 285 442 303
rect 507 309 509 319
rect 589 319 614 321
rect 529 306 531 311
rect 463 299 465 302
rect 462 297 468 299
rect 462 295 464 297
rect 466 295 468 297
rect 462 293 468 295
rect 440 274 442 277
rect 463 275 465 293
rect 473 289 475 303
rect 480 300 482 303
rect 480 298 486 300
rect 480 296 482 298
rect 484 296 486 298
rect 480 294 486 296
rect 490 290 492 303
rect 470 287 476 289
rect 470 285 472 287
rect 474 285 476 287
rect 470 283 476 285
rect 480 288 492 290
rect 497 294 499 303
rect 497 292 503 294
rect 497 290 499 292
rect 501 290 503 292
rect 497 288 503 290
rect 440 272 449 274
rect 443 270 445 272
rect 447 270 449 272
rect 443 268 449 270
rect 473 273 475 283
rect 480 273 482 288
rect 487 282 493 284
rect 487 280 489 282
rect 491 280 493 282
rect 487 278 493 280
rect 490 273 492 278
rect 497 273 499 288
rect 507 285 509 303
rect 539 303 541 308
rect 549 303 551 308
rect 572 314 574 319
rect 579 314 581 319
rect 589 311 591 319
rect 599 311 601 315
rect 612 311 614 319
rect 612 309 617 311
rect 615 306 617 309
rect 529 294 531 297
rect 539 294 541 297
rect 529 292 535 294
rect 529 290 531 292
rect 533 290 535 292
rect 529 288 535 290
rect 539 292 545 294
rect 539 290 541 292
rect 543 290 545 292
rect 539 288 545 290
rect 529 285 531 288
rect 507 274 509 277
rect 507 272 516 274
rect 510 270 512 272
rect 514 270 516 272
rect 510 268 516 270
rect 542 278 544 288
rect 549 287 551 297
rect 572 293 574 302
rect 579 299 581 302
rect 579 297 583 299
rect 589 298 591 302
rect 599 299 601 302
rect 581 294 583 297
rect 599 297 608 299
rect 599 295 604 297
rect 606 295 608 297
rect 571 291 577 293
rect 571 289 573 291
rect 575 289 577 291
rect 571 287 577 289
rect 581 292 587 294
rect 581 290 583 292
rect 585 290 587 292
rect 581 288 587 290
rect 599 293 608 295
rect 599 289 601 293
rect 615 289 617 297
rect 549 285 555 287
rect 549 283 551 285
rect 553 283 555 285
rect 571 284 573 287
rect 581 284 583 288
rect 591 287 601 289
rect 607 287 620 289
rect 591 284 593 287
rect 607 284 609 287
rect 618 286 620 287
rect 618 284 624 286
rect 549 281 555 283
rect 549 278 551 281
rect 529 262 531 267
rect 339 253 341 257
rect 346 253 348 257
rect 356 253 358 257
rect 363 253 365 257
rect 373 253 375 257
rect 396 253 398 257
rect 406 253 408 257
rect 413 253 415 257
rect 423 253 425 257
rect 430 253 432 257
rect 463 253 465 257
rect 473 253 475 257
rect 480 253 482 257
rect 490 253 492 257
rect 497 253 499 257
rect 581 262 583 266
rect 591 262 593 266
rect 542 253 544 257
rect 549 253 551 257
rect 571 253 573 257
rect 618 282 620 284
rect 622 282 624 284
rect 618 280 624 282
rect 607 253 609 257
rect 26 245 28 249
rect 33 245 35 249
rect 13 235 15 240
rect 110 245 112 249
rect 62 236 64 240
rect 72 238 74 243
rect 82 238 84 243
rect 13 214 15 217
rect 26 214 28 224
rect 33 221 35 224
rect 33 219 39 221
rect 33 217 35 219
rect 37 217 39 219
rect 33 215 39 217
rect 13 212 19 214
rect 13 210 15 212
rect 17 210 19 212
rect 13 208 19 210
rect 23 212 29 214
rect 23 210 25 212
rect 27 210 29 212
rect 23 208 29 210
rect 13 205 15 208
rect 23 205 25 208
rect 33 205 35 215
rect 62 214 64 218
rect 72 214 74 225
rect 82 222 84 225
rect 82 220 88 222
rect 82 218 84 220
rect 86 218 88 220
rect 82 216 88 218
rect 95 220 101 222
rect 95 218 97 220
rect 99 218 101 220
rect 146 245 148 249
rect 126 236 128 240
rect 136 236 138 240
rect 224 245 226 249
rect 176 236 178 240
rect 186 238 188 243
rect 196 238 198 243
rect 95 216 101 218
rect 62 212 68 214
rect 62 210 64 212
rect 66 210 68 212
rect 62 208 68 210
rect 72 212 78 214
rect 72 210 74 212
rect 76 210 78 212
rect 72 208 78 210
rect 62 203 64 208
rect 75 203 77 208
rect 82 203 84 216
rect 99 215 101 216
rect 110 215 112 218
rect 126 215 128 218
rect 99 213 112 215
rect 118 213 128 215
rect 136 214 138 218
rect 146 215 148 218
rect 102 205 104 213
rect 118 209 120 213
rect 111 207 120 209
rect 132 212 138 214
rect 132 210 134 212
rect 136 210 138 212
rect 132 208 138 210
rect 142 213 148 215
rect 142 211 144 213
rect 146 211 148 213
rect 142 209 148 211
rect 176 214 178 218
rect 186 214 188 225
rect 196 222 198 225
rect 196 220 202 222
rect 196 218 198 220
rect 200 218 202 220
rect 196 216 202 218
rect 209 220 215 222
rect 209 218 211 220
rect 213 218 215 220
rect 260 245 262 249
rect 240 236 242 240
rect 250 236 252 240
rect 339 245 341 249
rect 346 245 348 249
rect 356 245 358 249
rect 363 245 365 249
rect 373 245 375 249
rect 396 245 398 249
rect 406 245 408 249
rect 413 245 415 249
rect 423 245 425 249
rect 430 245 432 249
rect 463 245 465 249
rect 473 245 475 249
rect 480 245 482 249
rect 490 245 492 249
rect 497 245 499 249
rect 287 238 289 243
rect 297 238 299 243
rect 307 236 309 240
rect 287 222 289 225
rect 283 220 289 222
rect 283 218 285 220
rect 287 218 289 220
rect 209 216 215 218
rect 176 212 182 214
rect 176 210 178 212
rect 180 210 182 212
rect 111 205 113 207
rect 115 205 120 207
rect 13 191 15 196
rect 23 194 25 199
rect 33 194 35 199
rect 62 190 64 194
rect 111 203 120 205
rect 136 205 138 208
rect 118 200 120 203
rect 128 200 130 204
rect 136 203 140 205
rect 138 200 140 203
rect 145 200 147 209
rect 176 208 182 210
rect 186 212 192 214
rect 186 210 188 212
rect 190 210 192 212
rect 186 208 192 210
rect 176 203 178 208
rect 189 203 191 208
rect 196 203 198 216
rect 213 215 215 216
rect 224 215 226 218
rect 240 215 242 218
rect 213 213 226 215
rect 232 213 242 215
rect 250 214 252 218
rect 260 215 262 218
rect 283 216 289 218
rect 216 205 218 213
rect 232 209 234 213
rect 225 207 234 209
rect 246 212 252 214
rect 246 210 248 212
rect 250 210 252 212
rect 246 208 252 210
rect 256 213 262 215
rect 256 211 258 213
rect 260 211 262 213
rect 256 209 262 211
rect 225 205 227 207
rect 229 205 234 207
rect 102 193 104 196
rect 75 187 77 192
rect 82 187 84 192
rect 102 191 107 193
rect 105 183 107 191
rect 118 187 120 191
rect 128 183 130 191
rect 176 190 178 194
rect 225 203 234 205
rect 250 205 252 208
rect 232 200 234 203
rect 242 200 244 204
rect 250 203 254 205
rect 252 200 254 203
rect 259 200 261 209
rect 287 203 289 216
rect 297 214 299 225
rect 322 232 328 234
rect 322 230 324 232
rect 326 230 328 232
rect 322 228 331 230
rect 329 225 331 228
rect 307 214 309 218
rect 293 212 299 214
rect 293 210 295 212
rect 297 210 299 212
rect 293 208 299 210
rect 303 212 309 214
rect 303 210 305 212
rect 307 210 309 212
rect 303 208 309 210
rect 294 203 296 208
rect 307 203 309 208
rect 216 193 218 196
rect 138 183 140 188
rect 145 183 147 188
rect 105 181 130 183
rect 189 187 191 192
rect 196 187 198 192
rect 216 191 221 193
rect 219 183 221 191
rect 232 187 234 191
rect 242 183 244 191
rect 329 199 331 217
rect 339 214 341 229
rect 346 224 348 229
rect 345 222 351 224
rect 345 220 347 222
rect 349 220 351 222
rect 345 218 351 220
rect 356 214 358 229
rect 363 219 365 229
rect 443 232 449 234
rect 443 230 445 232
rect 447 230 449 232
rect 335 212 341 214
rect 335 210 337 212
rect 339 210 341 212
rect 335 208 341 210
rect 339 199 341 208
rect 346 212 358 214
rect 362 217 368 219
rect 362 215 364 217
rect 366 215 368 217
rect 362 213 368 215
rect 346 199 348 212
rect 352 206 358 208
rect 352 204 354 206
rect 356 204 358 206
rect 352 202 358 204
rect 356 199 358 202
rect 363 199 365 213
rect 373 209 375 227
rect 396 209 398 227
rect 406 219 408 229
rect 403 217 409 219
rect 403 215 405 217
rect 407 215 409 217
rect 403 213 409 215
rect 413 214 415 229
rect 423 224 425 229
rect 420 222 426 224
rect 420 220 422 222
rect 424 220 426 222
rect 420 218 426 220
rect 430 214 432 229
rect 440 228 449 230
rect 440 225 442 228
rect 542 245 544 249
rect 549 245 551 249
rect 571 245 573 249
rect 529 235 531 240
rect 510 232 516 234
rect 510 230 512 232
rect 514 230 516 232
rect 370 207 376 209
rect 370 205 372 207
rect 374 205 376 207
rect 370 203 376 205
rect 395 207 401 209
rect 395 205 397 207
rect 399 205 401 207
rect 395 203 401 205
rect 373 200 375 203
rect 396 200 398 203
rect 252 183 254 188
rect 259 183 261 188
rect 287 187 289 192
rect 294 187 296 192
rect 219 181 244 183
rect 307 190 309 194
rect 329 183 331 193
rect 406 199 408 213
rect 413 212 425 214
rect 413 206 419 208
rect 413 204 415 206
rect 417 204 419 206
rect 413 202 419 204
rect 413 199 415 202
rect 423 199 425 212
rect 430 212 436 214
rect 430 210 432 212
rect 434 210 436 212
rect 430 208 436 210
rect 430 199 432 208
rect 440 199 442 217
rect 463 209 465 227
rect 473 219 475 229
rect 470 217 476 219
rect 470 215 472 217
rect 474 215 476 217
rect 470 213 476 215
rect 480 214 482 229
rect 490 224 492 229
rect 487 222 493 224
rect 487 220 489 222
rect 491 220 493 222
rect 487 218 493 220
rect 497 214 499 229
rect 507 228 516 230
rect 507 225 509 228
rect 462 207 468 209
rect 462 205 464 207
rect 466 205 468 207
rect 462 203 468 205
rect 463 200 465 203
rect 339 187 341 191
rect 346 183 348 191
rect 356 186 358 191
rect 363 186 365 191
rect 373 186 375 191
rect 396 186 398 191
rect 406 186 408 191
rect 413 186 415 191
rect 329 181 348 183
rect 423 183 425 191
rect 430 187 432 191
rect 440 183 442 193
rect 473 199 475 213
rect 480 212 492 214
rect 480 206 486 208
rect 480 204 482 206
rect 484 204 486 206
rect 480 202 486 204
rect 480 199 482 202
rect 490 199 492 212
rect 497 212 503 214
rect 497 210 499 212
rect 501 210 503 212
rect 497 208 503 210
rect 497 199 499 208
rect 507 199 509 217
rect 529 214 531 217
rect 542 214 544 224
rect 549 221 551 224
rect 549 219 555 221
rect 549 217 551 219
rect 553 217 555 219
rect 607 245 609 249
rect 581 236 583 240
rect 591 236 593 240
rect 618 220 624 222
rect 618 218 620 220
rect 622 218 624 220
rect 549 215 555 217
rect 571 215 573 218
rect 529 212 535 214
rect 529 210 531 212
rect 533 210 535 212
rect 529 208 535 210
rect 539 212 545 214
rect 539 210 541 212
rect 543 210 545 212
rect 539 208 545 210
rect 529 205 531 208
rect 539 205 541 208
rect 549 205 551 215
rect 571 213 577 215
rect 571 211 573 213
rect 575 211 577 213
rect 571 209 577 211
rect 581 214 583 218
rect 591 215 593 218
rect 607 215 609 218
rect 618 216 624 218
rect 618 215 620 216
rect 581 212 587 214
rect 591 213 601 215
rect 607 213 620 215
rect 581 210 583 212
rect 585 210 587 212
rect 572 200 574 209
rect 581 208 587 210
rect 599 209 601 213
rect 581 205 583 208
rect 579 203 583 205
rect 599 207 608 209
rect 599 205 604 207
rect 606 205 608 207
rect 615 205 617 213
rect 579 200 581 203
rect 589 200 591 204
rect 599 203 608 205
rect 599 200 601 203
rect 463 186 465 191
rect 473 186 475 191
rect 480 186 482 191
rect 423 181 442 183
rect 490 183 492 191
rect 497 187 499 191
rect 507 183 509 193
rect 529 191 531 196
rect 539 194 541 199
rect 549 194 551 199
rect 490 181 509 183
rect 615 193 617 196
rect 612 191 617 193
rect 572 183 574 188
rect 579 183 581 188
rect 589 183 591 191
rect 599 187 601 191
rect 612 183 614 191
rect 589 181 614 183
rect 13 162 15 167
rect 23 159 25 164
rect 33 159 35 164
rect 62 164 64 168
rect 75 166 77 171
rect 82 166 84 171
rect 105 175 130 177
rect 105 167 107 175
rect 118 167 120 171
rect 128 167 130 175
rect 138 170 140 175
rect 145 170 147 175
rect 102 165 107 167
rect 102 162 104 165
rect 13 150 15 153
rect 23 150 25 153
rect 13 148 19 150
rect 13 146 15 148
rect 17 146 19 148
rect 13 144 19 146
rect 23 148 29 150
rect 23 146 25 148
rect 27 146 29 148
rect 23 144 29 146
rect 13 141 15 144
rect 26 134 28 144
rect 33 143 35 153
rect 62 150 64 155
rect 75 150 77 155
rect 62 148 68 150
rect 62 146 64 148
rect 66 146 68 148
rect 62 144 68 146
rect 72 148 78 150
rect 72 146 74 148
rect 76 146 78 148
rect 72 144 78 146
rect 33 141 39 143
rect 33 139 35 141
rect 37 139 39 141
rect 62 140 64 144
rect 33 137 39 139
rect 33 134 35 137
rect 13 118 15 123
rect 72 133 74 144
rect 82 142 84 155
rect 176 164 178 168
rect 189 166 191 171
rect 196 166 198 171
rect 219 175 244 177
rect 219 167 221 175
rect 232 167 234 171
rect 242 167 244 175
rect 252 170 254 175
rect 259 170 261 175
rect 118 155 120 158
rect 111 153 120 155
rect 128 154 130 158
rect 138 155 140 158
rect 102 145 104 153
rect 111 151 113 153
rect 115 151 120 153
rect 111 149 120 151
rect 136 153 140 155
rect 136 150 138 153
rect 118 145 120 149
rect 132 148 138 150
rect 145 149 147 158
rect 216 165 221 167
rect 216 162 218 165
rect 176 150 178 155
rect 189 150 191 155
rect 132 146 134 148
rect 136 146 138 148
rect 99 143 112 145
rect 118 143 128 145
rect 132 144 138 146
rect 99 142 101 143
rect 82 140 88 142
rect 82 138 84 140
rect 86 138 88 140
rect 82 136 88 138
rect 95 140 101 142
rect 110 140 112 143
rect 126 140 128 143
rect 136 140 138 144
rect 142 147 148 149
rect 142 145 144 147
rect 146 145 148 147
rect 142 143 148 145
rect 146 140 148 143
rect 176 148 182 150
rect 176 146 178 148
rect 180 146 182 148
rect 176 144 182 146
rect 186 148 192 150
rect 186 146 188 148
rect 190 146 192 148
rect 186 144 192 146
rect 176 140 178 144
rect 95 138 97 140
rect 99 138 101 140
rect 95 136 101 138
rect 82 133 84 136
rect 62 118 64 122
rect 72 115 74 120
rect 82 115 84 120
rect 26 109 28 113
rect 33 109 35 113
rect 126 118 128 122
rect 136 118 138 122
rect 110 109 112 113
rect 186 133 188 144
rect 196 142 198 155
rect 287 166 289 171
rect 294 166 296 171
rect 329 175 348 177
rect 232 155 234 158
rect 225 153 234 155
rect 242 154 244 158
rect 252 155 254 158
rect 216 145 218 153
rect 225 151 227 153
rect 229 151 234 153
rect 225 149 234 151
rect 250 153 254 155
rect 250 150 252 153
rect 232 145 234 149
rect 246 148 252 150
rect 259 149 261 158
rect 307 164 309 168
rect 329 165 331 175
rect 339 167 341 171
rect 346 167 348 175
rect 423 175 442 177
rect 356 167 358 172
rect 363 167 365 172
rect 373 167 375 172
rect 396 167 398 172
rect 406 167 408 172
rect 413 167 415 172
rect 423 167 425 175
rect 430 167 432 171
rect 246 146 248 148
rect 250 146 252 148
rect 213 143 226 145
rect 232 143 242 145
rect 246 144 252 146
rect 213 142 215 143
rect 196 140 202 142
rect 196 138 198 140
rect 200 138 202 140
rect 196 136 202 138
rect 209 140 215 142
rect 224 140 226 143
rect 240 140 242 143
rect 250 140 252 144
rect 256 147 262 149
rect 256 145 258 147
rect 260 145 262 147
rect 256 143 262 145
rect 260 140 262 143
rect 287 142 289 155
rect 294 150 296 155
rect 307 150 309 155
rect 293 148 299 150
rect 293 146 295 148
rect 297 146 299 148
rect 293 144 299 146
rect 303 148 309 150
rect 303 146 305 148
rect 307 146 309 148
rect 303 144 309 146
rect 283 140 289 142
rect 209 138 211 140
rect 213 138 215 140
rect 209 136 215 138
rect 196 133 198 136
rect 176 118 178 122
rect 186 115 188 120
rect 196 115 198 120
rect 146 109 148 113
rect 240 118 242 122
rect 250 118 252 122
rect 224 109 226 113
rect 283 138 285 140
rect 287 138 289 140
rect 283 136 289 138
rect 287 133 289 136
rect 297 133 299 144
rect 307 140 309 144
rect 329 141 331 159
rect 339 150 341 159
rect 335 148 341 150
rect 335 146 337 148
rect 339 146 341 148
rect 335 144 341 146
rect 346 146 348 159
rect 356 156 358 159
rect 352 154 358 156
rect 352 152 354 154
rect 356 152 358 154
rect 352 150 358 152
rect 346 144 358 146
rect 363 145 365 159
rect 440 165 442 175
rect 490 175 509 177
rect 463 167 465 172
rect 473 167 475 172
rect 480 167 482 172
rect 490 167 492 175
rect 497 167 499 171
rect 373 155 375 158
rect 396 155 398 158
rect 370 153 376 155
rect 370 151 372 153
rect 374 151 376 153
rect 370 149 376 151
rect 395 153 401 155
rect 395 151 397 153
rect 399 151 401 153
rect 395 149 401 151
rect 329 130 331 133
rect 322 128 331 130
rect 339 129 341 144
rect 345 138 351 140
rect 345 136 347 138
rect 349 136 351 138
rect 345 134 351 136
rect 346 129 348 134
rect 356 129 358 144
rect 362 143 368 145
rect 362 141 364 143
rect 366 141 368 143
rect 362 139 368 141
rect 363 129 365 139
rect 373 131 375 149
rect 396 131 398 149
rect 406 145 408 159
rect 413 156 415 159
rect 413 154 419 156
rect 413 152 415 154
rect 417 152 419 154
rect 413 150 419 152
rect 423 146 425 159
rect 403 143 409 145
rect 403 141 405 143
rect 407 141 409 143
rect 403 139 409 141
rect 413 144 425 146
rect 430 150 432 159
rect 430 148 436 150
rect 430 146 432 148
rect 434 146 436 148
rect 430 144 436 146
rect 322 126 324 128
rect 326 126 328 128
rect 322 124 328 126
rect 287 115 289 120
rect 297 115 299 120
rect 307 118 309 122
rect 260 109 262 113
rect 406 129 408 139
rect 413 129 415 144
rect 420 138 426 140
rect 420 136 422 138
rect 424 136 426 138
rect 420 134 426 136
rect 423 129 425 134
rect 430 129 432 144
rect 440 141 442 159
rect 507 165 509 175
rect 589 175 614 177
rect 529 162 531 167
rect 463 155 465 158
rect 462 153 468 155
rect 462 151 464 153
rect 466 151 468 153
rect 462 149 468 151
rect 440 130 442 133
rect 463 131 465 149
rect 473 145 475 159
rect 480 156 482 159
rect 480 154 486 156
rect 480 152 482 154
rect 484 152 486 154
rect 480 150 486 152
rect 490 146 492 159
rect 470 143 476 145
rect 470 141 472 143
rect 474 141 476 143
rect 470 139 476 141
rect 480 144 492 146
rect 497 150 499 159
rect 497 148 503 150
rect 497 146 499 148
rect 501 146 503 148
rect 497 144 503 146
rect 440 128 449 130
rect 443 126 445 128
rect 447 126 449 128
rect 443 124 449 126
rect 473 129 475 139
rect 480 129 482 144
rect 487 138 493 140
rect 487 136 489 138
rect 491 136 493 138
rect 487 134 493 136
rect 490 129 492 134
rect 497 129 499 144
rect 507 141 509 159
rect 539 159 541 164
rect 549 159 551 164
rect 572 170 574 175
rect 579 170 581 175
rect 589 167 591 175
rect 599 167 601 171
rect 612 167 614 175
rect 612 165 617 167
rect 615 162 617 165
rect 529 150 531 153
rect 539 150 541 153
rect 529 148 535 150
rect 529 146 531 148
rect 533 146 535 148
rect 529 144 535 146
rect 539 148 545 150
rect 539 146 541 148
rect 543 146 545 148
rect 539 144 545 146
rect 529 141 531 144
rect 507 130 509 133
rect 507 128 516 130
rect 510 126 512 128
rect 514 126 516 128
rect 510 124 516 126
rect 542 134 544 144
rect 549 143 551 153
rect 572 149 574 158
rect 579 155 581 158
rect 579 153 583 155
rect 589 154 591 158
rect 599 155 601 158
rect 581 150 583 153
rect 599 153 608 155
rect 599 151 604 153
rect 606 151 608 153
rect 571 147 577 149
rect 571 145 573 147
rect 575 145 577 147
rect 571 143 577 145
rect 581 148 587 150
rect 581 146 583 148
rect 585 146 587 148
rect 581 144 587 146
rect 599 149 608 151
rect 599 145 601 149
rect 615 145 617 153
rect 549 141 555 143
rect 549 139 551 141
rect 553 139 555 141
rect 571 140 573 143
rect 581 140 583 144
rect 591 143 601 145
rect 607 143 620 145
rect 591 140 593 143
rect 607 140 609 143
rect 618 142 620 143
rect 618 140 624 142
rect 549 137 555 139
rect 549 134 551 137
rect 529 118 531 123
rect 339 109 341 113
rect 346 109 348 113
rect 356 109 358 113
rect 363 109 365 113
rect 373 109 375 113
rect 396 109 398 113
rect 406 109 408 113
rect 413 109 415 113
rect 423 109 425 113
rect 430 109 432 113
rect 463 109 465 113
rect 473 109 475 113
rect 480 109 482 113
rect 490 109 492 113
rect 497 109 499 113
rect 581 118 583 122
rect 591 118 593 122
rect 542 109 544 113
rect 549 109 551 113
rect 571 109 573 113
rect 618 138 620 140
rect 622 138 624 140
rect 618 136 624 138
rect 607 109 609 113
rect 26 101 28 105
rect 33 101 35 105
rect 13 91 15 96
rect 110 101 112 105
rect 62 92 64 96
rect 72 94 74 99
rect 82 94 84 99
rect 13 70 15 73
rect 26 70 28 80
rect 33 77 35 80
rect 33 75 39 77
rect 33 73 35 75
rect 37 73 39 75
rect 33 71 39 73
rect 13 68 19 70
rect 13 66 15 68
rect 17 66 19 68
rect 13 64 19 66
rect 23 68 29 70
rect 23 66 25 68
rect 27 66 29 68
rect 23 64 29 66
rect 13 61 15 64
rect 23 61 25 64
rect 33 61 35 71
rect 62 70 64 74
rect 72 70 74 81
rect 82 78 84 81
rect 82 76 88 78
rect 82 74 84 76
rect 86 74 88 76
rect 82 72 88 74
rect 95 76 101 78
rect 95 74 97 76
rect 99 74 101 76
rect 146 101 148 105
rect 126 92 128 96
rect 136 92 138 96
rect 224 101 226 105
rect 176 92 178 96
rect 186 94 188 99
rect 196 94 198 99
rect 95 72 101 74
rect 62 68 68 70
rect 62 66 64 68
rect 66 66 68 68
rect 62 64 68 66
rect 72 68 78 70
rect 72 66 74 68
rect 76 66 78 68
rect 72 64 78 66
rect 62 59 64 64
rect 75 59 77 64
rect 82 59 84 72
rect 99 71 101 72
rect 110 71 112 74
rect 126 71 128 74
rect 99 69 112 71
rect 118 69 128 71
rect 136 70 138 74
rect 146 71 148 74
rect 102 61 104 69
rect 118 65 120 69
rect 111 63 120 65
rect 132 68 138 70
rect 132 66 134 68
rect 136 66 138 68
rect 132 64 138 66
rect 142 69 148 71
rect 142 67 144 69
rect 146 67 148 69
rect 142 65 148 67
rect 176 70 178 74
rect 186 70 188 81
rect 196 78 198 81
rect 196 76 202 78
rect 196 74 198 76
rect 200 74 202 76
rect 196 72 202 74
rect 209 76 215 78
rect 209 74 211 76
rect 213 74 215 76
rect 260 101 262 105
rect 240 92 242 96
rect 250 92 252 96
rect 339 101 341 105
rect 346 101 348 105
rect 356 101 358 105
rect 363 101 365 105
rect 373 101 375 105
rect 396 101 398 105
rect 406 101 408 105
rect 413 101 415 105
rect 423 101 425 105
rect 430 101 432 105
rect 463 101 465 105
rect 473 101 475 105
rect 480 101 482 105
rect 490 101 492 105
rect 497 101 499 105
rect 287 94 289 99
rect 297 94 299 99
rect 307 92 309 96
rect 287 78 289 81
rect 283 76 289 78
rect 283 74 285 76
rect 287 74 289 76
rect 209 72 215 74
rect 176 68 182 70
rect 176 66 178 68
rect 180 66 182 68
rect 111 61 113 63
rect 115 61 120 63
rect 13 47 15 52
rect 23 50 25 55
rect 33 50 35 55
rect 62 46 64 50
rect 111 59 120 61
rect 136 61 138 64
rect 118 56 120 59
rect 128 56 130 60
rect 136 59 140 61
rect 138 56 140 59
rect 145 56 147 65
rect 176 64 182 66
rect 186 68 192 70
rect 186 66 188 68
rect 190 66 192 68
rect 186 64 192 66
rect 176 59 178 64
rect 189 59 191 64
rect 196 59 198 72
rect 213 71 215 72
rect 224 71 226 74
rect 240 71 242 74
rect 213 69 226 71
rect 232 69 242 71
rect 250 70 252 74
rect 260 71 262 74
rect 283 72 289 74
rect 216 61 218 69
rect 232 65 234 69
rect 225 63 234 65
rect 246 68 252 70
rect 246 66 248 68
rect 250 66 252 68
rect 246 64 252 66
rect 256 69 262 71
rect 256 67 258 69
rect 260 67 262 69
rect 256 65 262 67
rect 225 61 227 63
rect 229 61 234 63
rect 102 49 104 52
rect 75 43 77 48
rect 82 43 84 48
rect 102 47 107 49
rect 105 39 107 47
rect 118 43 120 47
rect 128 39 130 47
rect 176 46 178 50
rect 225 59 234 61
rect 250 61 252 64
rect 232 56 234 59
rect 242 56 244 60
rect 250 59 254 61
rect 252 56 254 59
rect 259 56 261 65
rect 287 59 289 72
rect 297 70 299 81
rect 322 88 328 90
rect 322 86 324 88
rect 326 86 328 88
rect 322 84 331 86
rect 329 81 331 84
rect 307 70 309 74
rect 293 68 299 70
rect 293 66 295 68
rect 297 66 299 68
rect 293 64 299 66
rect 303 68 309 70
rect 303 66 305 68
rect 307 66 309 68
rect 303 64 309 66
rect 294 59 296 64
rect 307 59 309 64
rect 216 49 218 52
rect 138 39 140 44
rect 145 39 147 44
rect 105 37 130 39
rect 189 43 191 48
rect 196 43 198 48
rect 216 47 221 49
rect 219 39 221 47
rect 232 43 234 47
rect 242 39 244 47
rect 329 55 331 73
rect 339 70 341 85
rect 346 80 348 85
rect 345 78 351 80
rect 345 76 347 78
rect 349 76 351 78
rect 345 74 351 76
rect 356 70 358 85
rect 363 75 365 85
rect 443 88 449 90
rect 443 86 445 88
rect 447 86 449 88
rect 335 68 341 70
rect 335 66 337 68
rect 339 66 341 68
rect 335 64 341 66
rect 339 55 341 64
rect 346 68 358 70
rect 362 73 368 75
rect 362 71 364 73
rect 366 71 368 73
rect 362 69 368 71
rect 346 55 348 68
rect 352 62 358 64
rect 352 60 354 62
rect 356 60 358 62
rect 352 58 358 60
rect 356 55 358 58
rect 363 55 365 69
rect 373 65 375 83
rect 396 65 398 83
rect 406 75 408 85
rect 403 73 409 75
rect 403 71 405 73
rect 407 71 409 73
rect 403 69 409 71
rect 413 70 415 85
rect 423 80 425 85
rect 420 78 426 80
rect 420 76 422 78
rect 424 76 426 78
rect 420 74 426 76
rect 430 70 432 85
rect 440 84 449 86
rect 440 81 442 84
rect 542 101 544 105
rect 549 101 551 105
rect 571 101 573 105
rect 529 91 531 96
rect 510 88 516 90
rect 510 86 512 88
rect 514 86 516 88
rect 370 63 376 65
rect 370 61 372 63
rect 374 61 376 63
rect 370 59 376 61
rect 395 63 401 65
rect 395 61 397 63
rect 399 61 401 63
rect 395 59 401 61
rect 373 56 375 59
rect 396 56 398 59
rect 252 39 254 44
rect 259 39 261 44
rect 287 43 289 48
rect 294 43 296 48
rect 219 37 244 39
rect 307 46 309 50
rect 329 39 331 49
rect 406 55 408 69
rect 413 68 425 70
rect 413 62 419 64
rect 413 60 415 62
rect 417 60 419 62
rect 413 58 419 60
rect 413 55 415 58
rect 423 55 425 68
rect 430 68 436 70
rect 430 66 432 68
rect 434 66 436 68
rect 430 64 436 66
rect 430 55 432 64
rect 440 55 442 73
rect 463 65 465 83
rect 473 75 475 85
rect 470 73 476 75
rect 470 71 472 73
rect 474 71 476 73
rect 470 69 476 71
rect 480 70 482 85
rect 490 80 492 85
rect 487 78 493 80
rect 487 76 489 78
rect 491 76 493 78
rect 487 74 493 76
rect 497 70 499 85
rect 507 84 516 86
rect 507 81 509 84
rect 462 63 468 65
rect 462 61 464 63
rect 466 61 468 63
rect 462 59 468 61
rect 463 56 465 59
rect 339 43 341 47
rect 346 39 348 47
rect 356 42 358 47
rect 363 42 365 47
rect 373 42 375 47
rect 396 42 398 47
rect 406 42 408 47
rect 413 42 415 47
rect 329 37 348 39
rect 423 39 425 47
rect 430 43 432 47
rect 440 39 442 49
rect 473 55 475 69
rect 480 68 492 70
rect 480 62 486 64
rect 480 60 482 62
rect 484 60 486 62
rect 480 58 486 60
rect 480 55 482 58
rect 490 55 492 68
rect 497 68 503 70
rect 497 66 499 68
rect 501 66 503 68
rect 497 64 503 66
rect 497 55 499 64
rect 507 55 509 73
rect 529 70 531 73
rect 542 70 544 80
rect 549 77 551 80
rect 549 75 555 77
rect 549 73 551 75
rect 553 73 555 75
rect 607 101 609 105
rect 581 92 583 96
rect 591 92 593 96
rect 618 76 624 78
rect 618 74 620 76
rect 622 74 624 76
rect 549 71 555 73
rect 571 71 573 74
rect 529 68 535 70
rect 529 66 531 68
rect 533 66 535 68
rect 529 64 535 66
rect 539 68 545 70
rect 539 66 541 68
rect 543 66 545 68
rect 539 64 545 66
rect 529 61 531 64
rect 539 61 541 64
rect 549 61 551 71
rect 571 69 577 71
rect 571 67 573 69
rect 575 67 577 69
rect 571 65 577 67
rect 581 70 583 74
rect 591 71 593 74
rect 607 71 609 74
rect 618 72 624 74
rect 618 71 620 72
rect 581 68 587 70
rect 591 69 601 71
rect 607 69 620 71
rect 581 66 583 68
rect 585 66 587 68
rect 572 56 574 65
rect 581 64 587 66
rect 599 65 601 69
rect 581 61 583 64
rect 579 59 583 61
rect 599 63 608 65
rect 599 61 604 63
rect 606 61 608 63
rect 615 61 617 69
rect 579 56 581 59
rect 589 56 591 60
rect 599 59 608 61
rect 599 56 601 59
rect 463 42 465 47
rect 473 42 475 47
rect 480 42 482 47
rect 423 37 442 39
rect 490 39 492 47
rect 497 43 499 47
rect 507 39 509 49
rect 529 47 531 52
rect 539 50 541 55
rect 549 50 551 55
rect 490 37 509 39
rect 615 49 617 52
rect 612 47 617 49
rect 572 39 574 44
rect 579 39 581 44
rect 589 39 591 47
rect 599 43 601 47
rect 612 39 614 47
rect 589 37 614 39
<< ndif >>
rect 17 314 23 316
rect 17 312 19 314
rect 21 312 23 314
rect 17 310 23 312
rect 36 314 42 316
rect 66 318 73 320
rect 66 316 68 318
rect 70 316 73 318
rect 36 312 38 314
rect 40 312 42 314
rect 36 310 42 312
rect 17 306 21 310
rect 8 303 13 306
rect 6 301 13 303
rect 6 299 8 301
rect 10 299 13 301
rect 6 297 13 299
rect 15 303 21 306
rect 37 303 42 310
rect 66 310 73 316
rect 149 318 155 320
rect 149 316 151 318
rect 153 316 155 318
rect 149 314 155 316
rect 180 318 187 320
rect 180 316 182 318
rect 184 316 187 318
rect 133 311 138 314
rect 66 308 75 310
rect 15 297 23 303
rect 25 301 33 303
rect 25 299 28 301
rect 30 299 33 301
rect 25 297 33 299
rect 35 297 42 303
rect 55 306 62 308
rect 55 304 57 306
rect 59 304 62 306
rect 55 302 62 304
rect 57 299 62 302
rect 64 299 75 308
rect 77 299 82 310
rect 84 308 91 310
rect 84 306 87 308
rect 89 306 91 308
rect 109 309 118 311
rect 109 307 111 309
rect 113 307 118 309
rect 109 306 118 307
rect 84 304 91 306
rect 84 299 89 304
rect 97 303 102 306
rect 95 301 102 303
rect 95 299 97 301
rect 99 299 102 301
rect 95 297 102 299
rect 104 302 118 306
rect 120 306 128 311
rect 120 304 123 306
rect 125 304 128 306
rect 120 302 128 304
rect 130 308 138 311
rect 130 306 133 308
rect 135 306 138 308
rect 130 302 138 306
rect 140 302 145 314
rect 147 302 155 314
rect 180 310 187 316
rect 263 318 269 320
rect 263 316 265 318
rect 267 316 269 318
rect 263 314 269 316
rect 298 318 305 320
rect 298 316 301 318
rect 303 316 305 318
rect 247 311 252 314
rect 180 308 189 310
rect 169 306 176 308
rect 169 304 171 306
rect 173 304 176 306
rect 169 302 176 304
rect 104 297 109 302
rect 171 299 176 302
rect 178 299 189 308
rect 191 299 196 310
rect 198 308 205 310
rect 198 306 201 308
rect 203 306 205 308
rect 223 309 232 311
rect 223 307 225 309
rect 227 307 232 309
rect 223 306 232 307
rect 198 304 205 306
rect 198 299 203 304
rect 211 303 216 306
rect 209 301 216 303
rect 209 299 211 301
rect 213 299 216 301
rect 209 297 216 299
rect 218 302 232 306
rect 234 306 242 311
rect 234 304 237 306
rect 239 304 242 306
rect 234 302 242 304
rect 244 308 252 311
rect 244 306 247 308
rect 249 306 252 308
rect 244 302 252 306
rect 254 302 259 314
rect 261 302 269 314
rect 298 310 305 316
rect 280 308 287 310
rect 280 306 282 308
rect 284 306 287 308
rect 280 304 287 306
rect 218 297 223 302
rect 282 299 287 304
rect 289 299 294 310
rect 296 308 305 310
rect 333 309 339 311
rect 296 299 307 308
rect 309 306 316 308
rect 309 304 312 306
rect 314 304 316 306
rect 309 302 316 304
rect 322 307 329 309
rect 322 305 324 307
rect 326 305 329 307
rect 322 303 329 305
rect 331 307 339 309
rect 331 305 334 307
rect 336 305 339 307
rect 331 303 339 305
rect 341 303 346 311
rect 348 309 356 311
rect 348 307 351 309
rect 353 307 356 309
rect 348 303 356 307
rect 358 303 363 311
rect 365 309 373 311
rect 365 307 368 309
rect 370 307 373 309
rect 365 303 373 307
rect 309 299 314 302
rect 368 302 373 303
rect 375 308 380 311
rect 391 308 396 311
rect 375 306 382 308
rect 375 304 378 306
rect 380 304 382 306
rect 375 302 382 304
rect 389 306 396 308
rect 389 304 391 306
rect 393 304 396 306
rect 389 302 396 304
rect 398 309 406 311
rect 398 307 401 309
rect 403 307 406 309
rect 398 303 406 307
rect 408 303 413 311
rect 415 309 423 311
rect 415 307 418 309
rect 420 307 423 309
rect 415 303 423 307
rect 425 303 430 311
rect 432 309 438 311
rect 432 307 440 309
rect 432 305 435 307
rect 437 305 440 307
rect 432 303 440 305
rect 442 307 449 309
rect 458 308 463 311
rect 442 305 445 307
rect 447 305 449 307
rect 442 303 449 305
rect 456 306 463 308
rect 456 304 458 306
rect 460 304 463 306
rect 398 302 403 303
rect 456 302 463 304
rect 465 309 473 311
rect 465 307 468 309
rect 470 307 473 309
rect 465 303 473 307
rect 475 303 480 311
rect 482 309 490 311
rect 482 307 485 309
rect 487 307 490 309
rect 482 303 490 307
rect 492 303 497 311
rect 499 309 505 311
rect 564 318 570 320
rect 564 316 566 318
rect 568 316 570 318
rect 533 314 539 316
rect 533 312 535 314
rect 537 312 539 314
rect 499 307 507 309
rect 499 305 502 307
rect 504 305 507 307
rect 499 303 507 305
rect 509 307 516 309
rect 509 305 512 307
rect 514 305 516 307
rect 533 310 539 312
rect 552 314 558 316
rect 552 312 554 314
rect 556 312 558 314
rect 552 310 558 312
rect 533 306 537 310
rect 509 303 516 305
rect 524 303 529 306
rect 465 302 470 303
rect 522 301 529 303
rect 522 299 524 301
rect 526 299 529 301
rect 522 297 529 299
rect 531 303 537 306
rect 553 303 558 310
rect 531 297 539 303
rect 541 301 549 303
rect 541 299 544 301
rect 546 299 549 301
rect 541 297 549 299
rect 551 297 558 303
rect 564 314 570 316
rect 564 302 572 314
rect 574 302 579 314
rect 581 311 586 314
rect 581 308 589 311
rect 581 306 584 308
rect 586 306 589 308
rect 581 302 589 306
rect 591 306 599 311
rect 591 304 594 306
rect 596 304 599 306
rect 591 302 599 304
rect 601 309 610 311
rect 601 307 606 309
rect 608 307 610 309
rect 601 306 610 307
rect 601 302 615 306
rect 610 297 615 302
rect 617 303 622 306
rect 617 301 624 303
rect 617 299 620 301
rect 622 299 624 301
rect 617 297 624 299
rect 6 203 13 205
rect 6 201 8 203
rect 10 201 13 203
rect 6 199 13 201
rect 8 196 13 199
rect 15 199 23 205
rect 25 203 33 205
rect 25 201 28 203
rect 30 201 33 203
rect 25 199 33 201
rect 35 199 42 205
rect 95 203 102 205
rect 57 200 62 203
rect 15 196 21 199
rect 17 192 21 196
rect 37 192 42 199
rect 55 198 62 200
rect 55 196 57 198
rect 59 196 62 198
rect 55 194 62 196
rect 64 194 75 203
rect 17 190 23 192
rect 17 188 19 190
rect 21 188 23 190
rect 17 186 23 188
rect 36 190 42 192
rect 66 192 75 194
rect 77 192 82 203
rect 84 198 89 203
rect 95 201 97 203
rect 99 201 102 203
rect 95 199 102 201
rect 84 196 91 198
rect 97 196 102 199
rect 104 200 109 205
rect 209 203 216 205
rect 171 200 176 203
rect 104 196 118 200
rect 84 194 87 196
rect 89 194 91 196
rect 84 192 91 194
rect 109 195 118 196
rect 109 193 111 195
rect 113 193 118 195
rect 36 188 38 190
rect 40 188 42 190
rect 36 186 42 188
rect 66 186 73 192
rect 109 191 118 193
rect 120 198 128 200
rect 120 196 123 198
rect 125 196 128 198
rect 120 191 128 196
rect 130 196 138 200
rect 130 194 133 196
rect 135 194 138 196
rect 130 191 138 194
rect 66 184 68 186
rect 70 184 73 186
rect 66 182 73 184
rect 133 188 138 191
rect 140 188 145 200
rect 147 188 155 200
rect 169 198 176 200
rect 169 196 171 198
rect 173 196 176 198
rect 169 194 176 196
rect 178 194 189 203
rect 180 192 189 194
rect 191 192 196 203
rect 198 198 203 203
rect 209 201 211 203
rect 213 201 216 203
rect 209 199 216 201
rect 198 196 205 198
rect 211 196 216 199
rect 218 200 223 205
rect 218 196 232 200
rect 198 194 201 196
rect 203 194 205 196
rect 198 192 205 194
rect 223 195 232 196
rect 223 193 225 195
rect 227 193 232 195
rect 149 186 155 188
rect 149 184 151 186
rect 153 184 155 186
rect 149 182 155 184
rect 180 186 187 192
rect 223 191 232 193
rect 234 198 242 200
rect 234 196 237 198
rect 239 196 242 198
rect 234 191 242 196
rect 244 196 252 200
rect 244 194 247 196
rect 249 194 252 196
rect 244 191 252 194
rect 180 184 182 186
rect 184 184 187 186
rect 180 182 187 184
rect 247 188 252 191
rect 254 188 259 200
rect 261 188 269 200
rect 282 198 287 203
rect 280 196 287 198
rect 280 194 282 196
rect 284 194 287 196
rect 280 192 287 194
rect 289 192 294 203
rect 296 194 307 203
rect 309 200 314 203
rect 309 198 316 200
rect 368 199 373 200
rect 309 196 312 198
rect 314 196 316 198
rect 309 194 316 196
rect 322 197 329 199
rect 322 195 324 197
rect 326 195 329 197
rect 296 192 305 194
rect 263 186 269 188
rect 263 184 265 186
rect 267 184 269 186
rect 263 182 269 184
rect 298 186 305 192
rect 322 193 329 195
rect 331 197 339 199
rect 331 195 334 197
rect 336 195 339 197
rect 331 193 339 195
rect 298 184 301 186
rect 303 184 305 186
rect 298 182 305 184
rect 333 191 339 193
rect 341 191 346 199
rect 348 195 356 199
rect 348 193 351 195
rect 353 193 356 195
rect 348 191 356 193
rect 358 191 363 199
rect 365 195 373 199
rect 365 193 368 195
rect 370 193 373 195
rect 365 191 373 193
rect 375 198 382 200
rect 375 196 378 198
rect 380 196 382 198
rect 375 194 382 196
rect 389 198 396 200
rect 389 196 391 198
rect 393 196 396 198
rect 389 194 396 196
rect 375 191 380 194
rect 391 191 396 194
rect 398 199 403 200
rect 398 195 406 199
rect 398 193 401 195
rect 403 193 406 195
rect 398 191 406 193
rect 408 191 413 199
rect 415 195 423 199
rect 415 193 418 195
rect 420 193 423 195
rect 415 191 423 193
rect 425 191 430 199
rect 432 197 440 199
rect 432 195 435 197
rect 437 195 440 197
rect 432 193 440 195
rect 442 197 449 199
rect 442 195 445 197
rect 447 195 449 197
rect 442 193 449 195
rect 456 198 463 200
rect 456 196 458 198
rect 460 196 463 198
rect 456 194 463 196
rect 432 191 438 193
rect 458 191 463 194
rect 465 199 470 200
rect 522 203 529 205
rect 522 201 524 203
rect 526 201 529 203
rect 522 199 529 201
rect 465 195 473 199
rect 465 193 468 195
rect 470 193 473 195
rect 465 191 473 193
rect 475 191 480 199
rect 482 195 490 199
rect 482 193 485 195
rect 487 193 490 195
rect 482 191 490 193
rect 492 191 497 199
rect 499 197 507 199
rect 499 195 502 197
rect 504 195 507 197
rect 499 193 507 195
rect 509 197 516 199
rect 509 195 512 197
rect 514 195 516 197
rect 524 196 529 199
rect 531 199 539 205
rect 541 203 549 205
rect 541 201 544 203
rect 546 201 549 203
rect 541 199 549 201
rect 551 199 558 205
rect 610 200 615 205
rect 531 196 537 199
rect 509 193 516 195
rect 499 191 505 193
rect 533 192 537 196
rect 553 192 558 199
rect 533 190 539 192
rect 533 188 535 190
rect 537 188 539 190
rect 533 186 539 188
rect 552 190 558 192
rect 552 188 554 190
rect 556 188 558 190
rect 552 186 558 188
rect 564 188 572 200
rect 574 188 579 200
rect 581 196 589 200
rect 581 194 584 196
rect 586 194 589 196
rect 581 191 589 194
rect 591 198 599 200
rect 591 196 594 198
rect 596 196 599 198
rect 591 191 599 196
rect 601 196 615 200
rect 617 203 624 205
rect 617 201 620 203
rect 622 201 624 203
rect 617 199 624 201
rect 617 196 622 199
rect 601 195 610 196
rect 601 193 606 195
rect 608 193 610 195
rect 601 191 610 193
rect 581 188 586 191
rect 564 186 570 188
rect 564 184 566 186
rect 568 184 570 186
rect 564 182 570 184
rect 17 170 23 172
rect 17 168 19 170
rect 21 168 23 170
rect 17 166 23 168
rect 36 170 42 172
rect 66 174 73 176
rect 66 172 68 174
rect 70 172 73 174
rect 36 168 38 170
rect 40 168 42 170
rect 36 166 42 168
rect 17 162 21 166
rect 8 159 13 162
rect 6 157 13 159
rect 6 155 8 157
rect 10 155 13 157
rect 6 153 13 155
rect 15 159 21 162
rect 37 159 42 166
rect 66 166 73 172
rect 149 174 155 176
rect 149 172 151 174
rect 153 172 155 174
rect 149 170 155 172
rect 180 174 187 176
rect 180 172 182 174
rect 184 172 187 174
rect 133 167 138 170
rect 66 164 75 166
rect 15 153 23 159
rect 25 157 33 159
rect 25 155 28 157
rect 30 155 33 157
rect 25 153 33 155
rect 35 153 42 159
rect 55 162 62 164
rect 55 160 57 162
rect 59 160 62 162
rect 55 158 62 160
rect 57 155 62 158
rect 64 155 75 164
rect 77 155 82 166
rect 84 164 91 166
rect 84 162 87 164
rect 89 162 91 164
rect 109 165 118 167
rect 109 163 111 165
rect 113 163 118 165
rect 109 162 118 163
rect 84 160 91 162
rect 84 155 89 160
rect 97 159 102 162
rect 95 157 102 159
rect 95 155 97 157
rect 99 155 102 157
rect 95 153 102 155
rect 104 158 118 162
rect 120 162 128 167
rect 120 160 123 162
rect 125 160 128 162
rect 120 158 128 160
rect 130 164 138 167
rect 130 162 133 164
rect 135 162 138 164
rect 130 158 138 162
rect 140 158 145 170
rect 147 158 155 170
rect 180 166 187 172
rect 263 174 269 176
rect 263 172 265 174
rect 267 172 269 174
rect 263 170 269 172
rect 298 174 305 176
rect 298 172 301 174
rect 303 172 305 174
rect 247 167 252 170
rect 180 164 189 166
rect 169 162 176 164
rect 169 160 171 162
rect 173 160 176 162
rect 169 158 176 160
rect 104 153 109 158
rect 171 155 176 158
rect 178 155 189 164
rect 191 155 196 166
rect 198 164 205 166
rect 198 162 201 164
rect 203 162 205 164
rect 223 165 232 167
rect 223 163 225 165
rect 227 163 232 165
rect 223 162 232 163
rect 198 160 205 162
rect 198 155 203 160
rect 211 159 216 162
rect 209 157 216 159
rect 209 155 211 157
rect 213 155 216 157
rect 209 153 216 155
rect 218 158 232 162
rect 234 162 242 167
rect 234 160 237 162
rect 239 160 242 162
rect 234 158 242 160
rect 244 164 252 167
rect 244 162 247 164
rect 249 162 252 164
rect 244 158 252 162
rect 254 158 259 170
rect 261 158 269 170
rect 298 166 305 172
rect 280 164 287 166
rect 280 162 282 164
rect 284 162 287 164
rect 280 160 287 162
rect 218 153 223 158
rect 282 155 287 160
rect 289 155 294 166
rect 296 164 305 166
rect 333 165 339 167
rect 296 155 307 164
rect 309 162 316 164
rect 309 160 312 162
rect 314 160 316 162
rect 309 158 316 160
rect 322 163 329 165
rect 322 161 324 163
rect 326 161 329 163
rect 322 159 329 161
rect 331 163 339 165
rect 331 161 334 163
rect 336 161 339 163
rect 331 159 339 161
rect 341 159 346 167
rect 348 165 356 167
rect 348 163 351 165
rect 353 163 356 165
rect 348 159 356 163
rect 358 159 363 167
rect 365 165 373 167
rect 365 163 368 165
rect 370 163 373 165
rect 365 159 373 163
rect 309 155 314 158
rect 368 158 373 159
rect 375 164 380 167
rect 391 164 396 167
rect 375 162 382 164
rect 375 160 378 162
rect 380 160 382 162
rect 375 158 382 160
rect 389 162 396 164
rect 389 160 391 162
rect 393 160 396 162
rect 389 158 396 160
rect 398 165 406 167
rect 398 163 401 165
rect 403 163 406 165
rect 398 159 406 163
rect 408 159 413 167
rect 415 165 423 167
rect 415 163 418 165
rect 420 163 423 165
rect 415 159 423 163
rect 425 159 430 167
rect 432 165 438 167
rect 432 163 440 165
rect 432 161 435 163
rect 437 161 440 163
rect 432 159 440 161
rect 442 163 449 165
rect 458 164 463 167
rect 442 161 445 163
rect 447 161 449 163
rect 442 159 449 161
rect 456 162 463 164
rect 456 160 458 162
rect 460 160 463 162
rect 398 158 403 159
rect 456 158 463 160
rect 465 165 473 167
rect 465 163 468 165
rect 470 163 473 165
rect 465 159 473 163
rect 475 159 480 167
rect 482 165 490 167
rect 482 163 485 165
rect 487 163 490 165
rect 482 159 490 163
rect 492 159 497 167
rect 499 165 505 167
rect 564 174 570 176
rect 564 172 566 174
rect 568 172 570 174
rect 533 170 539 172
rect 533 168 535 170
rect 537 168 539 170
rect 499 163 507 165
rect 499 161 502 163
rect 504 161 507 163
rect 499 159 507 161
rect 509 163 516 165
rect 509 161 512 163
rect 514 161 516 163
rect 533 166 539 168
rect 552 170 558 172
rect 552 168 554 170
rect 556 168 558 170
rect 552 166 558 168
rect 533 162 537 166
rect 509 159 516 161
rect 524 159 529 162
rect 465 158 470 159
rect 522 157 529 159
rect 522 155 524 157
rect 526 155 529 157
rect 522 153 529 155
rect 531 159 537 162
rect 553 159 558 166
rect 531 153 539 159
rect 541 157 549 159
rect 541 155 544 157
rect 546 155 549 157
rect 541 153 549 155
rect 551 153 558 159
rect 564 170 570 172
rect 564 158 572 170
rect 574 158 579 170
rect 581 167 586 170
rect 581 164 589 167
rect 581 162 584 164
rect 586 162 589 164
rect 581 158 589 162
rect 591 162 599 167
rect 591 160 594 162
rect 596 160 599 162
rect 591 158 599 160
rect 601 165 610 167
rect 601 163 606 165
rect 608 163 610 165
rect 601 162 610 163
rect 601 158 615 162
rect 610 153 615 158
rect 617 159 622 162
rect 617 157 624 159
rect 617 155 620 157
rect 622 155 624 157
rect 617 153 624 155
rect 6 59 13 61
rect 6 57 8 59
rect 10 57 13 59
rect 6 55 13 57
rect 8 52 13 55
rect 15 55 23 61
rect 25 59 33 61
rect 25 57 28 59
rect 30 57 33 59
rect 25 55 33 57
rect 35 55 42 61
rect 95 59 102 61
rect 57 56 62 59
rect 15 52 21 55
rect 17 48 21 52
rect 37 48 42 55
rect 55 54 62 56
rect 55 52 57 54
rect 59 52 62 54
rect 55 50 62 52
rect 64 50 75 59
rect 17 46 23 48
rect 17 44 19 46
rect 21 44 23 46
rect 17 42 23 44
rect 36 46 42 48
rect 66 48 75 50
rect 77 48 82 59
rect 84 54 89 59
rect 95 57 97 59
rect 99 57 102 59
rect 95 55 102 57
rect 84 52 91 54
rect 97 52 102 55
rect 104 56 109 61
rect 209 59 216 61
rect 171 56 176 59
rect 104 52 118 56
rect 84 50 87 52
rect 89 50 91 52
rect 84 48 91 50
rect 109 51 118 52
rect 109 49 111 51
rect 113 49 118 51
rect 36 44 38 46
rect 40 44 42 46
rect 36 42 42 44
rect 66 42 73 48
rect 109 47 118 49
rect 120 54 128 56
rect 120 52 123 54
rect 125 52 128 54
rect 120 47 128 52
rect 130 52 138 56
rect 130 50 133 52
rect 135 50 138 52
rect 130 47 138 50
rect 66 40 68 42
rect 70 40 73 42
rect 66 38 73 40
rect 133 44 138 47
rect 140 44 145 56
rect 147 44 155 56
rect 169 54 176 56
rect 169 52 171 54
rect 173 52 176 54
rect 169 50 176 52
rect 178 50 189 59
rect 180 48 189 50
rect 191 48 196 59
rect 198 54 203 59
rect 209 57 211 59
rect 213 57 216 59
rect 209 55 216 57
rect 198 52 205 54
rect 211 52 216 55
rect 218 56 223 61
rect 218 52 232 56
rect 198 50 201 52
rect 203 50 205 52
rect 198 48 205 50
rect 223 51 232 52
rect 223 49 225 51
rect 227 49 232 51
rect 149 42 155 44
rect 149 40 151 42
rect 153 40 155 42
rect 149 38 155 40
rect 180 42 187 48
rect 223 47 232 49
rect 234 54 242 56
rect 234 52 237 54
rect 239 52 242 54
rect 234 47 242 52
rect 244 52 252 56
rect 244 50 247 52
rect 249 50 252 52
rect 244 47 252 50
rect 180 40 182 42
rect 184 40 187 42
rect 180 38 187 40
rect 247 44 252 47
rect 254 44 259 56
rect 261 44 269 56
rect 282 54 287 59
rect 280 52 287 54
rect 280 50 282 52
rect 284 50 287 52
rect 280 48 287 50
rect 289 48 294 59
rect 296 50 307 59
rect 309 56 314 59
rect 309 54 316 56
rect 368 55 373 56
rect 309 52 312 54
rect 314 52 316 54
rect 309 50 316 52
rect 322 53 329 55
rect 322 51 324 53
rect 326 51 329 53
rect 296 48 305 50
rect 263 42 269 44
rect 263 40 265 42
rect 267 40 269 42
rect 263 38 269 40
rect 298 42 305 48
rect 322 49 329 51
rect 331 53 339 55
rect 331 51 334 53
rect 336 51 339 53
rect 331 49 339 51
rect 298 40 301 42
rect 303 40 305 42
rect 298 38 305 40
rect 333 47 339 49
rect 341 47 346 55
rect 348 51 356 55
rect 348 49 351 51
rect 353 49 356 51
rect 348 47 356 49
rect 358 47 363 55
rect 365 51 373 55
rect 365 49 368 51
rect 370 49 373 51
rect 365 47 373 49
rect 375 54 382 56
rect 375 52 378 54
rect 380 52 382 54
rect 375 50 382 52
rect 389 54 396 56
rect 389 52 391 54
rect 393 52 396 54
rect 389 50 396 52
rect 375 47 380 50
rect 391 47 396 50
rect 398 55 403 56
rect 398 51 406 55
rect 398 49 401 51
rect 403 49 406 51
rect 398 47 406 49
rect 408 47 413 55
rect 415 51 423 55
rect 415 49 418 51
rect 420 49 423 51
rect 415 47 423 49
rect 425 47 430 55
rect 432 53 440 55
rect 432 51 435 53
rect 437 51 440 53
rect 432 49 440 51
rect 442 53 449 55
rect 442 51 445 53
rect 447 51 449 53
rect 442 49 449 51
rect 456 54 463 56
rect 456 52 458 54
rect 460 52 463 54
rect 456 50 463 52
rect 432 47 438 49
rect 458 47 463 50
rect 465 55 470 56
rect 522 59 529 61
rect 522 57 524 59
rect 526 57 529 59
rect 522 55 529 57
rect 465 51 473 55
rect 465 49 468 51
rect 470 49 473 51
rect 465 47 473 49
rect 475 47 480 55
rect 482 51 490 55
rect 482 49 485 51
rect 487 49 490 51
rect 482 47 490 49
rect 492 47 497 55
rect 499 53 507 55
rect 499 51 502 53
rect 504 51 507 53
rect 499 49 507 51
rect 509 53 516 55
rect 509 51 512 53
rect 514 51 516 53
rect 524 52 529 55
rect 531 55 539 61
rect 541 59 549 61
rect 541 57 544 59
rect 546 57 549 59
rect 541 55 549 57
rect 551 55 558 61
rect 610 56 615 61
rect 531 52 537 55
rect 509 49 516 51
rect 499 47 505 49
rect 533 48 537 52
rect 553 48 558 55
rect 533 46 539 48
rect 533 44 535 46
rect 537 44 539 46
rect 533 42 539 44
rect 552 46 558 48
rect 552 44 554 46
rect 556 44 558 46
rect 552 42 558 44
rect 564 44 572 56
rect 574 44 579 56
rect 581 52 589 56
rect 581 50 584 52
rect 586 50 589 52
rect 581 47 589 50
rect 591 54 599 56
rect 591 52 594 54
rect 596 52 599 54
rect 591 47 599 52
rect 601 52 615 56
rect 617 59 624 61
rect 617 57 620 59
rect 622 57 624 59
rect 617 55 624 57
rect 617 52 622 55
rect 601 51 610 52
rect 601 49 606 51
rect 608 49 610 51
rect 601 47 610 49
rect 581 44 586 47
rect 564 42 570 44
rect 564 40 566 42
rect 568 40 570 42
rect 564 38 570 40
<< pdif >>
rect 8 280 13 285
rect 6 278 13 280
rect 6 276 8 278
rect 10 276 13 278
rect 6 271 13 276
rect 6 269 8 271
rect 10 269 13 271
rect 6 267 13 269
rect 15 278 23 285
rect 55 282 62 284
rect 55 280 57 282
rect 59 280 62 282
rect 15 267 26 278
rect 17 261 26 267
rect 17 259 19 261
rect 21 259 26 261
rect 17 257 26 259
rect 28 257 33 278
rect 35 270 40 278
rect 55 275 62 280
rect 55 273 57 275
rect 59 273 62 275
rect 55 271 62 273
rect 35 268 42 270
rect 35 266 38 268
rect 40 266 42 268
rect 57 266 62 271
rect 64 277 70 284
rect 103 282 110 284
rect 103 280 105 282
rect 107 280 110 282
rect 103 278 110 280
rect 64 270 72 277
rect 64 268 67 270
rect 69 268 72 270
rect 64 266 72 268
rect 35 264 42 266
rect 35 257 40 264
rect 66 264 72 266
rect 74 275 82 277
rect 74 273 77 275
rect 79 273 82 275
rect 74 268 82 273
rect 74 266 77 268
rect 79 266 82 268
rect 74 264 82 266
rect 84 268 91 277
rect 84 266 87 268
rect 89 266 91 268
rect 84 264 91 266
rect 105 257 110 278
rect 112 268 126 284
rect 112 266 115 268
rect 117 266 126 268
rect 128 282 136 284
rect 128 280 131 282
rect 133 280 136 282
rect 128 275 136 280
rect 128 273 131 275
rect 133 273 136 275
rect 128 266 136 273
rect 138 275 146 284
rect 138 273 141 275
rect 143 273 146 275
rect 138 266 146 273
rect 112 261 124 266
rect 112 259 115 261
rect 117 259 124 261
rect 112 257 124 259
rect 141 257 146 266
rect 148 269 153 284
rect 169 282 176 284
rect 169 280 171 282
rect 173 280 176 282
rect 169 275 176 280
rect 169 273 171 275
rect 173 273 176 275
rect 169 271 176 273
rect 148 267 155 269
rect 148 265 151 267
rect 153 265 155 267
rect 171 266 176 271
rect 178 277 184 284
rect 217 282 224 284
rect 217 280 219 282
rect 221 280 224 282
rect 217 278 224 280
rect 178 270 186 277
rect 178 268 181 270
rect 183 268 186 270
rect 178 266 186 268
rect 148 263 155 265
rect 148 257 153 263
rect 180 264 186 266
rect 188 275 196 277
rect 188 273 191 275
rect 193 273 196 275
rect 188 268 196 273
rect 188 266 191 268
rect 193 266 196 268
rect 188 264 196 266
rect 198 268 205 277
rect 198 266 201 268
rect 203 266 205 268
rect 198 264 205 266
rect 219 257 224 278
rect 226 268 240 284
rect 226 266 229 268
rect 231 266 240 268
rect 242 282 250 284
rect 242 280 245 282
rect 247 280 250 282
rect 242 275 250 280
rect 242 273 245 275
rect 247 273 250 275
rect 242 266 250 273
rect 252 275 260 284
rect 252 273 255 275
rect 257 273 260 275
rect 252 266 260 273
rect 226 261 238 266
rect 226 259 229 261
rect 231 259 238 261
rect 226 257 238 259
rect 255 257 260 266
rect 262 269 267 284
rect 301 277 307 284
rect 262 267 269 269
rect 262 265 265 267
rect 267 265 269 267
rect 262 263 269 265
rect 280 268 287 277
rect 280 266 282 268
rect 284 266 287 268
rect 280 264 287 266
rect 289 275 297 277
rect 289 273 292 275
rect 294 273 297 275
rect 289 268 297 273
rect 289 266 292 268
rect 294 266 297 268
rect 289 264 297 266
rect 299 270 307 277
rect 299 268 302 270
rect 304 268 307 270
rect 299 266 307 268
rect 309 282 316 284
rect 309 280 312 282
rect 314 280 316 282
rect 309 275 316 280
rect 322 283 329 285
rect 322 281 324 283
rect 326 281 329 283
rect 322 279 329 281
rect 324 277 329 279
rect 331 277 337 285
rect 309 273 312 275
rect 314 273 316 275
rect 309 271 316 273
rect 333 273 337 277
rect 368 273 373 275
rect 309 266 314 271
rect 333 269 339 273
rect 299 264 305 266
rect 262 257 267 263
rect 332 261 339 269
rect 332 259 334 261
rect 336 259 339 261
rect 332 257 339 259
rect 341 257 346 273
rect 348 271 356 273
rect 348 269 351 271
rect 353 269 356 271
rect 348 257 356 269
rect 358 257 363 273
rect 365 261 373 273
rect 365 259 368 261
rect 370 259 373 261
rect 365 257 373 259
rect 375 270 380 275
rect 391 270 396 275
rect 375 268 382 270
rect 375 266 378 268
rect 380 266 382 268
rect 375 264 382 266
rect 389 268 396 270
rect 389 266 391 268
rect 393 266 396 268
rect 389 264 396 266
rect 375 257 380 264
rect 391 257 396 264
rect 398 273 403 275
rect 434 277 440 285
rect 442 283 449 285
rect 442 281 445 283
rect 447 281 449 283
rect 442 279 449 281
rect 442 277 447 279
rect 434 273 438 277
rect 398 261 406 273
rect 398 259 401 261
rect 403 259 406 261
rect 398 257 406 259
rect 408 257 413 273
rect 415 271 423 273
rect 415 269 418 271
rect 420 269 423 271
rect 415 257 423 269
rect 425 257 430 273
rect 432 269 438 273
rect 458 270 463 275
rect 432 261 439 269
rect 456 268 463 270
rect 456 266 458 268
rect 460 266 463 268
rect 456 264 463 266
rect 432 259 435 261
rect 437 259 439 261
rect 432 257 439 259
rect 458 257 463 264
rect 465 273 470 275
rect 501 277 507 285
rect 509 283 516 285
rect 509 281 512 283
rect 514 281 516 283
rect 509 279 516 281
rect 524 280 529 285
rect 509 277 514 279
rect 522 278 529 280
rect 501 273 505 277
rect 465 261 473 273
rect 465 259 468 261
rect 470 259 473 261
rect 465 257 473 259
rect 475 257 480 273
rect 482 271 490 273
rect 482 269 485 271
rect 487 269 490 271
rect 482 257 490 269
rect 492 257 497 273
rect 499 269 505 273
rect 522 276 524 278
rect 526 276 529 278
rect 499 261 506 269
rect 522 271 529 276
rect 522 269 524 271
rect 526 269 529 271
rect 522 267 529 269
rect 531 278 539 285
rect 531 267 542 278
rect 499 259 502 261
rect 504 259 506 261
rect 533 261 542 267
rect 499 257 506 259
rect 533 259 535 261
rect 537 259 542 261
rect 533 257 542 259
rect 544 257 549 278
rect 551 270 556 278
rect 551 268 558 270
rect 566 269 571 284
rect 551 266 554 268
rect 556 266 558 268
rect 551 264 558 266
rect 564 267 571 269
rect 564 265 566 267
rect 568 265 571 267
rect 551 257 556 264
rect 564 263 571 265
rect 566 257 571 263
rect 573 275 581 284
rect 573 273 576 275
rect 578 273 581 275
rect 573 266 581 273
rect 583 282 591 284
rect 583 280 586 282
rect 588 280 591 282
rect 583 275 591 280
rect 583 273 586 275
rect 588 273 591 275
rect 583 266 591 273
rect 593 268 607 284
rect 593 266 602 268
rect 604 266 607 268
rect 573 257 578 266
rect 595 261 607 266
rect 595 259 602 261
rect 604 259 607 261
rect 595 257 607 259
rect 609 282 616 284
rect 609 280 612 282
rect 614 280 616 282
rect 609 278 616 280
rect 609 257 614 278
rect 17 243 26 245
rect 17 241 19 243
rect 21 241 26 243
rect 17 235 26 241
rect 6 233 13 235
rect 6 231 8 233
rect 10 231 13 233
rect 6 226 13 231
rect 6 224 8 226
rect 10 224 13 226
rect 6 222 13 224
rect 8 217 13 222
rect 15 224 26 235
rect 28 224 33 245
rect 35 238 40 245
rect 35 236 42 238
rect 66 236 72 238
rect 35 234 38 236
rect 40 234 42 236
rect 35 232 42 234
rect 35 224 40 232
rect 57 231 62 236
rect 55 229 62 231
rect 55 227 57 229
rect 59 227 62 229
rect 15 217 23 224
rect 55 222 62 227
rect 55 220 57 222
rect 59 220 62 222
rect 55 218 62 220
rect 64 234 72 236
rect 64 232 67 234
rect 69 232 72 234
rect 64 225 72 232
rect 74 236 82 238
rect 74 234 77 236
rect 79 234 82 236
rect 74 229 82 234
rect 74 227 77 229
rect 79 227 82 229
rect 74 225 82 227
rect 84 236 91 238
rect 84 234 87 236
rect 89 234 91 236
rect 84 225 91 234
rect 64 218 70 225
rect 105 224 110 245
rect 103 222 110 224
rect 103 220 105 222
rect 107 220 110 222
rect 103 218 110 220
rect 112 243 124 245
rect 112 241 115 243
rect 117 241 124 243
rect 112 236 124 241
rect 141 236 146 245
rect 112 234 115 236
rect 117 234 126 236
rect 112 218 126 234
rect 128 229 136 236
rect 128 227 131 229
rect 133 227 136 229
rect 128 222 136 227
rect 128 220 131 222
rect 133 220 136 222
rect 128 218 136 220
rect 138 229 146 236
rect 138 227 141 229
rect 143 227 146 229
rect 138 218 146 227
rect 148 239 153 245
rect 148 237 155 239
rect 148 235 151 237
rect 153 235 155 237
rect 180 236 186 238
rect 148 233 155 235
rect 148 218 153 233
rect 171 231 176 236
rect 169 229 176 231
rect 169 227 171 229
rect 173 227 176 229
rect 169 222 176 227
rect 169 220 171 222
rect 173 220 176 222
rect 169 218 176 220
rect 178 234 186 236
rect 178 232 181 234
rect 183 232 186 234
rect 178 225 186 232
rect 188 236 196 238
rect 188 234 191 236
rect 193 234 196 236
rect 188 229 196 234
rect 188 227 191 229
rect 193 227 196 229
rect 188 225 196 227
rect 198 236 205 238
rect 198 234 201 236
rect 203 234 205 236
rect 198 225 205 234
rect 178 218 184 225
rect 219 224 224 245
rect 217 222 224 224
rect 217 220 219 222
rect 221 220 224 222
rect 217 218 224 220
rect 226 243 238 245
rect 226 241 229 243
rect 231 241 238 243
rect 226 236 238 241
rect 255 236 260 245
rect 226 234 229 236
rect 231 234 240 236
rect 226 218 240 234
rect 242 229 250 236
rect 242 227 245 229
rect 247 227 250 229
rect 242 222 250 227
rect 242 220 245 222
rect 247 220 250 222
rect 242 218 250 220
rect 252 229 260 236
rect 252 227 255 229
rect 257 227 260 229
rect 252 218 260 227
rect 262 239 267 245
rect 262 237 269 239
rect 332 243 339 245
rect 332 241 334 243
rect 336 241 339 243
rect 262 235 265 237
rect 267 235 269 237
rect 262 233 269 235
rect 280 236 287 238
rect 280 234 282 236
rect 284 234 287 236
rect 262 218 267 233
rect 280 225 287 234
rect 289 236 297 238
rect 289 234 292 236
rect 294 234 297 236
rect 289 229 297 234
rect 289 227 292 229
rect 294 227 297 229
rect 289 225 297 227
rect 299 236 305 238
rect 299 234 307 236
rect 299 232 302 234
rect 304 232 307 234
rect 299 225 307 232
rect 301 218 307 225
rect 309 231 314 236
rect 332 233 339 241
rect 309 229 316 231
rect 309 227 312 229
rect 314 227 316 229
rect 309 222 316 227
rect 333 229 339 233
rect 341 229 346 245
rect 348 233 356 245
rect 348 231 351 233
rect 353 231 356 233
rect 348 229 356 231
rect 358 229 363 245
rect 365 243 373 245
rect 365 241 368 243
rect 370 241 373 243
rect 365 229 373 241
rect 333 225 337 229
rect 324 223 329 225
rect 309 220 312 222
rect 314 220 316 222
rect 309 218 316 220
rect 322 221 329 223
rect 322 219 324 221
rect 326 219 329 221
rect 322 217 329 219
rect 331 217 337 225
rect 368 227 373 229
rect 375 238 380 245
rect 391 238 396 245
rect 375 236 382 238
rect 375 234 378 236
rect 380 234 382 236
rect 375 232 382 234
rect 389 236 396 238
rect 389 234 391 236
rect 393 234 396 236
rect 389 232 396 234
rect 375 227 380 232
rect 391 227 396 232
rect 398 243 406 245
rect 398 241 401 243
rect 403 241 406 243
rect 398 229 406 241
rect 408 229 413 245
rect 415 233 423 245
rect 415 231 418 233
rect 420 231 423 233
rect 415 229 423 231
rect 425 229 430 245
rect 432 243 439 245
rect 432 241 435 243
rect 437 241 439 243
rect 432 233 439 241
rect 458 238 463 245
rect 456 236 463 238
rect 456 234 458 236
rect 460 234 463 236
rect 432 229 438 233
rect 456 232 463 234
rect 398 227 403 229
rect 434 225 438 229
rect 458 227 463 232
rect 465 243 473 245
rect 465 241 468 243
rect 470 241 473 243
rect 465 229 473 241
rect 475 229 480 245
rect 482 233 490 245
rect 482 231 485 233
rect 487 231 490 233
rect 482 229 490 231
rect 492 229 497 245
rect 499 243 506 245
rect 499 241 502 243
rect 504 241 506 243
rect 533 243 542 245
rect 499 233 506 241
rect 533 241 535 243
rect 537 241 542 243
rect 533 235 542 241
rect 499 229 505 233
rect 465 227 470 229
rect 434 217 440 225
rect 442 223 447 225
rect 442 221 449 223
rect 442 219 445 221
rect 447 219 449 221
rect 442 217 449 219
rect 501 225 505 229
rect 522 233 529 235
rect 522 231 524 233
rect 526 231 529 233
rect 522 226 529 231
rect 501 217 507 225
rect 509 223 514 225
rect 522 224 524 226
rect 526 224 529 226
rect 509 221 516 223
rect 522 222 529 224
rect 509 219 512 221
rect 514 219 516 221
rect 509 217 516 219
rect 524 217 529 222
rect 531 224 542 235
rect 544 224 549 245
rect 551 238 556 245
rect 566 239 571 245
rect 551 236 558 238
rect 551 234 554 236
rect 556 234 558 236
rect 551 232 558 234
rect 564 237 571 239
rect 564 235 566 237
rect 568 235 571 237
rect 564 233 571 235
rect 551 224 556 232
rect 531 217 539 224
rect 566 218 571 233
rect 573 236 578 245
rect 595 243 607 245
rect 595 241 602 243
rect 604 241 607 243
rect 595 236 607 241
rect 573 229 581 236
rect 573 227 576 229
rect 578 227 581 229
rect 573 218 581 227
rect 583 229 591 236
rect 583 227 586 229
rect 588 227 591 229
rect 583 222 591 227
rect 583 220 586 222
rect 588 220 591 222
rect 583 218 591 220
rect 593 234 602 236
rect 604 234 607 236
rect 593 218 607 234
rect 609 224 614 245
rect 609 222 616 224
rect 609 220 612 222
rect 614 220 616 222
rect 609 218 616 220
rect 8 136 13 141
rect 6 134 13 136
rect 6 132 8 134
rect 10 132 13 134
rect 6 127 13 132
rect 6 125 8 127
rect 10 125 13 127
rect 6 123 13 125
rect 15 134 23 141
rect 55 138 62 140
rect 55 136 57 138
rect 59 136 62 138
rect 15 123 26 134
rect 17 117 26 123
rect 17 115 19 117
rect 21 115 26 117
rect 17 113 26 115
rect 28 113 33 134
rect 35 126 40 134
rect 55 131 62 136
rect 55 129 57 131
rect 59 129 62 131
rect 55 127 62 129
rect 35 124 42 126
rect 35 122 38 124
rect 40 122 42 124
rect 57 122 62 127
rect 64 133 70 140
rect 103 138 110 140
rect 103 136 105 138
rect 107 136 110 138
rect 103 134 110 136
rect 64 126 72 133
rect 64 124 67 126
rect 69 124 72 126
rect 64 122 72 124
rect 35 120 42 122
rect 35 113 40 120
rect 66 120 72 122
rect 74 131 82 133
rect 74 129 77 131
rect 79 129 82 131
rect 74 124 82 129
rect 74 122 77 124
rect 79 122 82 124
rect 74 120 82 122
rect 84 124 91 133
rect 84 122 87 124
rect 89 122 91 124
rect 84 120 91 122
rect 105 113 110 134
rect 112 124 126 140
rect 112 122 115 124
rect 117 122 126 124
rect 128 138 136 140
rect 128 136 131 138
rect 133 136 136 138
rect 128 131 136 136
rect 128 129 131 131
rect 133 129 136 131
rect 128 122 136 129
rect 138 131 146 140
rect 138 129 141 131
rect 143 129 146 131
rect 138 122 146 129
rect 112 117 124 122
rect 112 115 115 117
rect 117 115 124 117
rect 112 113 124 115
rect 141 113 146 122
rect 148 125 153 140
rect 169 138 176 140
rect 169 136 171 138
rect 173 136 176 138
rect 169 131 176 136
rect 169 129 171 131
rect 173 129 176 131
rect 169 127 176 129
rect 148 123 155 125
rect 148 121 151 123
rect 153 121 155 123
rect 171 122 176 127
rect 178 133 184 140
rect 217 138 224 140
rect 217 136 219 138
rect 221 136 224 138
rect 217 134 224 136
rect 178 126 186 133
rect 178 124 181 126
rect 183 124 186 126
rect 178 122 186 124
rect 148 119 155 121
rect 148 113 153 119
rect 180 120 186 122
rect 188 131 196 133
rect 188 129 191 131
rect 193 129 196 131
rect 188 124 196 129
rect 188 122 191 124
rect 193 122 196 124
rect 188 120 196 122
rect 198 124 205 133
rect 198 122 201 124
rect 203 122 205 124
rect 198 120 205 122
rect 219 113 224 134
rect 226 124 240 140
rect 226 122 229 124
rect 231 122 240 124
rect 242 138 250 140
rect 242 136 245 138
rect 247 136 250 138
rect 242 131 250 136
rect 242 129 245 131
rect 247 129 250 131
rect 242 122 250 129
rect 252 131 260 140
rect 252 129 255 131
rect 257 129 260 131
rect 252 122 260 129
rect 226 117 238 122
rect 226 115 229 117
rect 231 115 238 117
rect 226 113 238 115
rect 255 113 260 122
rect 262 125 267 140
rect 301 133 307 140
rect 262 123 269 125
rect 262 121 265 123
rect 267 121 269 123
rect 262 119 269 121
rect 280 124 287 133
rect 280 122 282 124
rect 284 122 287 124
rect 280 120 287 122
rect 289 131 297 133
rect 289 129 292 131
rect 294 129 297 131
rect 289 124 297 129
rect 289 122 292 124
rect 294 122 297 124
rect 289 120 297 122
rect 299 126 307 133
rect 299 124 302 126
rect 304 124 307 126
rect 299 122 307 124
rect 309 138 316 140
rect 309 136 312 138
rect 314 136 316 138
rect 309 131 316 136
rect 322 139 329 141
rect 322 137 324 139
rect 326 137 329 139
rect 322 135 329 137
rect 324 133 329 135
rect 331 133 337 141
rect 309 129 312 131
rect 314 129 316 131
rect 309 127 316 129
rect 333 129 337 133
rect 368 129 373 131
rect 309 122 314 127
rect 333 125 339 129
rect 299 120 305 122
rect 262 113 267 119
rect 332 117 339 125
rect 332 115 334 117
rect 336 115 339 117
rect 332 113 339 115
rect 341 113 346 129
rect 348 127 356 129
rect 348 125 351 127
rect 353 125 356 127
rect 348 113 356 125
rect 358 113 363 129
rect 365 117 373 129
rect 365 115 368 117
rect 370 115 373 117
rect 365 113 373 115
rect 375 126 380 131
rect 391 126 396 131
rect 375 124 382 126
rect 375 122 378 124
rect 380 122 382 124
rect 375 120 382 122
rect 389 124 396 126
rect 389 122 391 124
rect 393 122 396 124
rect 389 120 396 122
rect 375 113 380 120
rect 391 113 396 120
rect 398 129 403 131
rect 434 133 440 141
rect 442 139 449 141
rect 442 137 445 139
rect 447 137 449 139
rect 442 135 449 137
rect 442 133 447 135
rect 434 129 438 133
rect 398 117 406 129
rect 398 115 401 117
rect 403 115 406 117
rect 398 113 406 115
rect 408 113 413 129
rect 415 127 423 129
rect 415 125 418 127
rect 420 125 423 127
rect 415 113 423 125
rect 425 113 430 129
rect 432 125 438 129
rect 458 126 463 131
rect 432 117 439 125
rect 456 124 463 126
rect 456 122 458 124
rect 460 122 463 124
rect 456 120 463 122
rect 432 115 435 117
rect 437 115 439 117
rect 432 113 439 115
rect 458 113 463 120
rect 465 129 470 131
rect 501 133 507 141
rect 509 139 516 141
rect 509 137 512 139
rect 514 137 516 139
rect 509 135 516 137
rect 524 136 529 141
rect 509 133 514 135
rect 522 134 529 136
rect 501 129 505 133
rect 465 117 473 129
rect 465 115 468 117
rect 470 115 473 117
rect 465 113 473 115
rect 475 113 480 129
rect 482 127 490 129
rect 482 125 485 127
rect 487 125 490 127
rect 482 113 490 125
rect 492 113 497 129
rect 499 125 505 129
rect 522 132 524 134
rect 526 132 529 134
rect 499 117 506 125
rect 522 127 529 132
rect 522 125 524 127
rect 526 125 529 127
rect 522 123 529 125
rect 531 134 539 141
rect 531 123 542 134
rect 499 115 502 117
rect 504 115 506 117
rect 533 117 542 123
rect 499 113 506 115
rect 533 115 535 117
rect 537 115 542 117
rect 533 113 542 115
rect 544 113 549 134
rect 551 126 556 134
rect 551 124 558 126
rect 566 125 571 140
rect 551 122 554 124
rect 556 122 558 124
rect 551 120 558 122
rect 564 123 571 125
rect 564 121 566 123
rect 568 121 571 123
rect 551 113 556 120
rect 564 119 571 121
rect 566 113 571 119
rect 573 131 581 140
rect 573 129 576 131
rect 578 129 581 131
rect 573 122 581 129
rect 583 138 591 140
rect 583 136 586 138
rect 588 136 591 138
rect 583 131 591 136
rect 583 129 586 131
rect 588 129 591 131
rect 583 122 591 129
rect 593 124 607 140
rect 593 122 602 124
rect 604 122 607 124
rect 573 113 578 122
rect 595 117 607 122
rect 595 115 602 117
rect 604 115 607 117
rect 595 113 607 115
rect 609 138 616 140
rect 609 136 612 138
rect 614 136 616 138
rect 609 134 616 136
rect 609 113 614 134
rect 17 99 26 101
rect 17 97 19 99
rect 21 97 26 99
rect 17 91 26 97
rect 6 89 13 91
rect 6 87 8 89
rect 10 87 13 89
rect 6 82 13 87
rect 6 80 8 82
rect 10 80 13 82
rect 6 78 13 80
rect 8 73 13 78
rect 15 80 26 91
rect 28 80 33 101
rect 35 94 40 101
rect 35 92 42 94
rect 66 92 72 94
rect 35 90 38 92
rect 40 90 42 92
rect 35 88 42 90
rect 35 80 40 88
rect 57 87 62 92
rect 55 85 62 87
rect 55 83 57 85
rect 59 83 62 85
rect 15 73 23 80
rect 55 78 62 83
rect 55 76 57 78
rect 59 76 62 78
rect 55 74 62 76
rect 64 90 72 92
rect 64 88 67 90
rect 69 88 72 90
rect 64 81 72 88
rect 74 92 82 94
rect 74 90 77 92
rect 79 90 82 92
rect 74 85 82 90
rect 74 83 77 85
rect 79 83 82 85
rect 74 81 82 83
rect 84 92 91 94
rect 84 90 87 92
rect 89 90 91 92
rect 84 81 91 90
rect 64 74 70 81
rect 105 80 110 101
rect 103 78 110 80
rect 103 76 105 78
rect 107 76 110 78
rect 103 74 110 76
rect 112 99 124 101
rect 112 97 115 99
rect 117 97 124 99
rect 112 92 124 97
rect 141 92 146 101
rect 112 90 115 92
rect 117 90 126 92
rect 112 74 126 90
rect 128 85 136 92
rect 128 83 131 85
rect 133 83 136 85
rect 128 78 136 83
rect 128 76 131 78
rect 133 76 136 78
rect 128 74 136 76
rect 138 85 146 92
rect 138 83 141 85
rect 143 83 146 85
rect 138 74 146 83
rect 148 95 153 101
rect 148 93 155 95
rect 148 91 151 93
rect 153 91 155 93
rect 180 92 186 94
rect 148 89 155 91
rect 148 74 153 89
rect 171 87 176 92
rect 169 85 176 87
rect 169 83 171 85
rect 173 83 176 85
rect 169 78 176 83
rect 169 76 171 78
rect 173 76 176 78
rect 169 74 176 76
rect 178 90 186 92
rect 178 88 181 90
rect 183 88 186 90
rect 178 81 186 88
rect 188 92 196 94
rect 188 90 191 92
rect 193 90 196 92
rect 188 85 196 90
rect 188 83 191 85
rect 193 83 196 85
rect 188 81 196 83
rect 198 92 205 94
rect 198 90 201 92
rect 203 90 205 92
rect 198 81 205 90
rect 178 74 184 81
rect 219 80 224 101
rect 217 78 224 80
rect 217 76 219 78
rect 221 76 224 78
rect 217 74 224 76
rect 226 99 238 101
rect 226 97 229 99
rect 231 97 238 99
rect 226 92 238 97
rect 255 92 260 101
rect 226 90 229 92
rect 231 90 240 92
rect 226 74 240 90
rect 242 85 250 92
rect 242 83 245 85
rect 247 83 250 85
rect 242 78 250 83
rect 242 76 245 78
rect 247 76 250 78
rect 242 74 250 76
rect 252 85 260 92
rect 252 83 255 85
rect 257 83 260 85
rect 252 74 260 83
rect 262 95 267 101
rect 262 93 269 95
rect 332 99 339 101
rect 332 97 334 99
rect 336 97 339 99
rect 262 91 265 93
rect 267 91 269 93
rect 262 89 269 91
rect 280 92 287 94
rect 280 90 282 92
rect 284 90 287 92
rect 262 74 267 89
rect 280 81 287 90
rect 289 92 297 94
rect 289 90 292 92
rect 294 90 297 92
rect 289 85 297 90
rect 289 83 292 85
rect 294 83 297 85
rect 289 81 297 83
rect 299 92 305 94
rect 299 90 307 92
rect 299 88 302 90
rect 304 88 307 90
rect 299 81 307 88
rect 301 74 307 81
rect 309 87 314 92
rect 332 89 339 97
rect 309 85 316 87
rect 309 83 312 85
rect 314 83 316 85
rect 309 78 316 83
rect 333 85 339 89
rect 341 85 346 101
rect 348 89 356 101
rect 348 87 351 89
rect 353 87 356 89
rect 348 85 356 87
rect 358 85 363 101
rect 365 99 373 101
rect 365 97 368 99
rect 370 97 373 99
rect 365 85 373 97
rect 333 81 337 85
rect 324 79 329 81
rect 309 76 312 78
rect 314 76 316 78
rect 309 74 316 76
rect 322 77 329 79
rect 322 75 324 77
rect 326 75 329 77
rect 322 73 329 75
rect 331 73 337 81
rect 368 83 373 85
rect 375 94 380 101
rect 391 94 396 101
rect 375 92 382 94
rect 375 90 378 92
rect 380 90 382 92
rect 375 88 382 90
rect 389 92 396 94
rect 389 90 391 92
rect 393 90 396 92
rect 389 88 396 90
rect 375 83 380 88
rect 391 83 396 88
rect 398 99 406 101
rect 398 97 401 99
rect 403 97 406 99
rect 398 85 406 97
rect 408 85 413 101
rect 415 89 423 101
rect 415 87 418 89
rect 420 87 423 89
rect 415 85 423 87
rect 425 85 430 101
rect 432 99 439 101
rect 432 97 435 99
rect 437 97 439 99
rect 432 89 439 97
rect 458 94 463 101
rect 456 92 463 94
rect 456 90 458 92
rect 460 90 463 92
rect 432 85 438 89
rect 456 88 463 90
rect 398 83 403 85
rect 434 81 438 85
rect 458 83 463 88
rect 465 99 473 101
rect 465 97 468 99
rect 470 97 473 99
rect 465 85 473 97
rect 475 85 480 101
rect 482 89 490 101
rect 482 87 485 89
rect 487 87 490 89
rect 482 85 490 87
rect 492 85 497 101
rect 499 99 506 101
rect 499 97 502 99
rect 504 97 506 99
rect 533 99 542 101
rect 499 89 506 97
rect 533 97 535 99
rect 537 97 542 99
rect 533 91 542 97
rect 499 85 505 89
rect 465 83 470 85
rect 434 73 440 81
rect 442 79 447 81
rect 442 77 449 79
rect 442 75 445 77
rect 447 75 449 77
rect 442 73 449 75
rect 501 81 505 85
rect 522 89 529 91
rect 522 87 524 89
rect 526 87 529 89
rect 522 82 529 87
rect 501 73 507 81
rect 509 79 514 81
rect 522 80 524 82
rect 526 80 529 82
rect 509 77 516 79
rect 522 78 529 80
rect 509 75 512 77
rect 514 75 516 77
rect 509 73 516 75
rect 524 73 529 78
rect 531 80 542 91
rect 544 80 549 101
rect 551 94 556 101
rect 566 95 571 101
rect 551 92 558 94
rect 551 90 554 92
rect 556 90 558 92
rect 551 88 558 90
rect 564 93 571 95
rect 564 91 566 93
rect 568 91 571 93
rect 564 89 571 91
rect 551 80 556 88
rect 531 73 539 80
rect 566 74 571 89
rect 573 92 578 101
rect 595 99 607 101
rect 595 97 602 99
rect 604 97 607 99
rect 595 92 607 97
rect 573 85 581 92
rect 573 83 576 85
rect 578 83 581 85
rect 573 74 581 83
rect 583 85 591 92
rect 583 83 586 85
rect 588 83 591 85
rect 583 78 591 83
rect 583 76 586 78
rect 588 76 591 78
rect 583 74 591 76
rect 593 90 602 92
rect 604 90 607 92
rect 593 74 607 90
rect 609 80 614 101
rect 609 78 616 80
rect 609 76 612 78
rect 614 76 616 78
rect 609 74 616 76
<< alu1 >>
rect 2 318 632 323
rect 2 316 9 318
rect 11 316 58 318
rect 60 316 68 318
rect 70 316 98 318
rect 100 316 151 318
rect 153 316 172 318
rect 174 316 182 318
rect 184 316 212 318
rect 214 316 265 318
rect 267 316 301 318
rect 303 316 311 318
rect 313 316 525 318
rect 527 316 566 318
rect 568 316 619 318
rect 621 316 632 318
rect 2 315 632 316
rect 55 306 67 310
rect 55 304 57 306
rect 59 304 67 306
rect 131 308 155 309
rect 6 301 11 303
rect 6 299 8 301
rect 10 299 11 301
rect 6 297 11 299
rect 6 278 10 297
rect 38 293 42 302
rect 6 276 8 278
rect 6 271 10 276
rect 6 269 8 271
rect 21 292 42 293
rect 21 290 25 292
rect 27 290 39 292
rect 41 290 42 292
rect 21 289 42 290
rect 21 283 35 285
rect 37 283 42 285
rect 21 281 42 283
rect 38 279 42 281
rect 55 284 59 304
rect 131 306 133 308
rect 135 306 155 308
rect 131 305 155 306
rect 79 301 84 302
rect 79 299 80 301
rect 82 299 84 301
rect 79 293 84 299
rect 55 282 60 284
rect 55 280 57 282
rect 59 280 60 282
rect 55 279 60 280
rect 38 275 60 279
rect 38 272 42 275
rect 55 273 57 275
rect 59 273 60 275
rect 70 292 84 293
rect 70 290 74 292
rect 76 290 84 292
rect 70 289 84 290
rect 103 301 116 302
rect 103 299 105 301
rect 107 299 116 301
rect 103 297 116 299
rect 103 296 113 297
rect 111 295 113 296
rect 115 295 116 297
rect 78 284 91 285
rect 78 282 84 284
rect 86 282 91 284
rect 78 281 91 282
rect 55 271 60 273
rect 6 265 19 269
rect 6 264 10 265
rect 87 277 91 281
rect 87 275 88 277
rect 90 275 91 277
rect 87 272 91 275
rect 95 284 100 286
rect 95 282 97 284
rect 99 282 100 284
rect 95 277 100 282
rect 111 288 116 295
rect 151 300 155 305
rect 151 298 152 300
rect 154 298 155 300
rect 95 275 97 277
rect 99 275 100 277
rect 95 270 100 275
rect 95 264 107 270
rect 151 277 155 298
rect 139 275 155 277
rect 139 273 141 275
rect 143 273 155 275
rect 139 272 155 273
rect 169 306 181 310
rect 169 304 171 306
rect 173 304 181 306
rect 245 308 269 309
rect 169 292 173 304
rect 245 306 247 308
rect 249 306 269 308
rect 245 305 269 306
rect 169 290 170 292
rect 172 290 173 292
rect 169 284 173 290
rect 193 301 198 302
rect 193 299 194 301
rect 196 299 198 301
rect 193 293 198 299
rect 169 282 174 284
rect 169 280 171 282
rect 173 280 174 282
rect 169 275 174 280
rect 169 273 171 275
rect 173 273 174 275
rect 184 292 198 293
rect 184 290 188 292
rect 190 290 198 292
rect 184 289 198 290
rect 217 301 230 302
rect 217 299 219 301
rect 221 299 230 301
rect 217 297 230 299
rect 217 296 227 297
rect 225 295 227 296
rect 229 295 230 297
rect 192 284 205 285
rect 192 282 198 284
rect 200 282 205 284
rect 192 281 205 282
rect 169 271 174 273
rect 201 277 205 281
rect 201 275 202 277
rect 204 275 205 277
rect 201 272 205 275
rect 209 284 214 286
rect 209 282 211 284
rect 213 282 214 284
rect 209 277 214 282
rect 225 288 230 295
rect 209 275 211 277
rect 213 275 214 277
rect 209 270 214 275
rect 209 264 221 270
rect 265 285 269 305
rect 287 293 292 302
rect 304 306 316 310
rect 304 304 312 306
rect 314 304 316 306
rect 287 292 301 293
rect 287 290 295 292
rect 297 290 301 292
rect 287 289 301 290
rect 265 283 266 285
rect 268 283 269 285
rect 265 277 269 283
rect 253 275 269 277
rect 253 273 255 275
rect 257 273 269 275
rect 253 272 269 273
rect 280 284 293 285
rect 280 282 285 284
rect 287 282 293 284
rect 280 281 293 282
rect 280 272 284 281
rect 312 300 316 304
rect 312 298 313 300
rect 315 298 316 300
rect 312 284 316 298
rect 311 282 316 284
rect 311 280 312 282
rect 314 280 316 282
rect 378 308 382 310
rect 377 306 382 308
rect 377 304 378 306
rect 380 304 382 306
rect 377 302 382 304
rect 329 300 342 301
rect 329 298 330 300
rect 332 298 342 300
rect 329 297 342 298
rect 336 292 342 297
rect 336 290 337 292
rect 339 290 342 292
rect 336 288 342 290
rect 362 287 366 294
rect 362 286 364 287
rect 354 285 364 286
rect 354 284 366 285
rect 354 282 355 284
rect 357 282 366 284
rect 354 280 366 282
rect 311 275 316 280
rect 311 273 312 275
rect 314 273 316 275
rect 311 271 316 273
rect 322 276 335 277
rect 322 274 332 276
rect 334 274 335 276
rect 322 273 335 274
rect 322 272 327 273
rect 378 292 382 302
rect 378 290 379 292
rect 381 290 382 292
rect 322 270 324 272
rect 326 270 327 272
rect 322 264 327 270
rect 378 269 382 290
rect 369 268 382 269
rect 369 266 378 268
rect 380 266 382 268
rect 369 265 382 266
rect 389 308 393 310
rect 389 306 394 308
rect 389 304 391 306
rect 393 304 394 306
rect 456 308 460 310
rect 389 302 394 304
rect 389 269 393 302
rect 429 300 442 301
rect 405 292 409 294
rect 405 290 406 292
rect 408 290 409 292
rect 405 287 409 290
rect 407 286 409 287
rect 407 285 417 286
rect 405 280 417 285
rect 429 298 437 300
rect 439 298 442 300
rect 429 297 442 298
rect 429 292 435 297
rect 429 290 432 292
rect 434 290 435 292
rect 429 288 435 290
rect 456 306 461 308
rect 456 304 458 306
rect 460 304 461 306
rect 564 308 588 309
rect 456 302 461 304
rect 456 300 460 302
rect 456 298 457 300
rect 459 298 460 300
rect 496 300 509 301
rect 436 273 449 277
rect 444 272 449 273
rect 389 268 402 269
rect 444 270 445 272
rect 447 270 449 272
rect 389 266 391 268
rect 393 266 402 268
rect 389 265 402 266
rect 444 264 449 270
rect 456 269 460 298
rect 472 287 476 294
rect 474 286 476 287
rect 474 285 484 286
rect 472 283 480 285
rect 482 283 484 285
rect 472 280 484 283
rect 496 298 505 300
rect 507 298 509 300
rect 496 297 509 298
rect 496 292 502 297
rect 496 290 499 292
rect 501 290 502 292
rect 496 288 502 290
rect 564 306 584 308
rect 586 306 588 308
rect 564 305 588 306
rect 522 301 527 303
rect 522 299 524 301
rect 526 299 527 301
rect 522 297 527 299
rect 522 284 526 297
rect 522 282 523 284
rect 525 282 526 284
rect 522 278 526 282
rect 554 293 558 302
rect 503 276 516 277
rect 503 274 504 276
rect 506 274 516 276
rect 503 273 516 274
rect 511 272 516 273
rect 456 268 469 269
rect 511 270 512 272
rect 514 270 516 272
rect 456 266 458 268
rect 460 266 469 268
rect 456 265 469 266
rect 511 264 516 270
rect 522 276 524 278
rect 522 271 526 276
rect 522 269 524 271
rect 537 292 558 293
rect 537 290 541 292
rect 543 290 558 292
rect 537 289 558 290
rect 564 300 568 305
rect 564 298 565 300
rect 567 298 568 300
rect 537 283 551 285
rect 553 283 558 285
rect 537 281 558 283
rect 554 272 558 281
rect 564 277 568 298
rect 603 297 616 302
rect 603 295 604 297
rect 606 296 616 297
rect 606 295 608 296
rect 564 275 580 277
rect 564 273 576 275
rect 578 273 580 275
rect 564 272 580 273
rect 603 288 608 295
rect 619 284 624 286
rect 619 282 620 284
rect 622 282 624 284
rect 522 265 535 269
rect 619 270 624 282
rect 522 264 526 265
rect 612 264 624 270
rect 2 258 632 259
rect 2 256 9 258
rect 11 256 58 258
rect 60 256 131 258
rect 133 256 172 258
rect 174 256 245 258
rect 247 256 311 258
rect 313 256 525 258
rect 527 256 586 258
rect 588 256 632 258
rect 2 246 632 256
rect 2 244 9 246
rect 11 244 58 246
rect 60 244 131 246
rect 133 244 172 246
rect 174 244 245 246
rect 247 244 311 246
rect 313 244 525 246
rect 527 244 586 246
rect 588 244 632 246
rect 2 243 632 244
rect 6 237 10 238
rect 6 233 19 237
rect 6 231 8 233
rect 6 226 10 231
rect 6 224 8 226
rect 6 221 10 224
rect 38 227 42 230
rect 55 229 60 231
rect 55 227 57 229
rect 59 227 60 229
rect 95 232 107 238
rect 6 219 7 221
rect 9 219 10 221
rect 6 205 10 219
rect 38 223 60 227
rect 38 221 42 223
rect 21 219 42 221
rect 21 217 35 219
rect 37 217 42 219
rect 55 222 60 223
rect 55 220 57 222
rect 59 220 60 222
rect 55 218 60 220
rect 87 227 91 230
rect 87 225 88 227
rect 90 225 91 227
rect 6 203 11 205
rect 6 201 8 203
rect 10 201 11 203
rect 6 199 11 201
rect 21 212 42 213
rect 21 210 25 212
rect 27 210 39 212
rect 41 210 42 212
rect 21 209 42 210
rect 38 200 42 209
rect 55 198 59 218
rect 87 221 91 225
rect 78 220 91 221
rect 78 218 84 220
rect 86 218 91 220
rect 78 217 91 218
rect 95 227 100 232
rect 95 225 97 227
rect 99 225 100 227
rect 95 220 100 225
rect 95 218 97 220
rect 99 218 100 220
rect 95 216 100 218
rect 70 212 84 213
rect 70 210 74 212
rect 76 210 84 212
rect 70 209 84 210
rect 55 196 57 198
rect 59 196 67 198
rect 55 192 67 196
rect 79 203 84 209
rect 79 201 80 203
rect 82 201 84 203
rect 79 200 84 201
rect 111 207 116 214
rect 139 229 155 230
rect 139 227 141 229
rect 143 227 155 229
rect 139 225 155 227
rect 111 206 113 207
rect 103 205 113 206
rect 115 205 116 207
rect 103 203 116 205
rect 103 201 105 203
rect 107 201 116 203
rect 103 200 116 201
rect 151 204 155 225
rect 151 202 152 204
rect 154 202 155 204
rect 151 197 155 202
rect 131 196 155 197
rect 131 194 133 196
rect 135 194 155 196
rect 131 193 155 194
rect 169 229 174 231
rect 169 227 171 229
rect 173 227 174 229
rect 209 232 221 238
rect 169 222 174 227
rect 169 220 171 222
rect 173 220 174 222
rect 169 218 174 220
rect 201 227 205 230
rect 201 225 202 227
rect 204 225 205 227
rect 169 212 173 218
rect 169 210 170 212
rect 172 210 173 212
rect 169 198 173 210
rect 201 221 205 225
rect 192 220 205 221
rect 192 218 198 220
rect 200 218 205 220
rect 192 217 205 218
rect 209 227 214 232
rect 209 225 211 227
rect 213 225 214 227
rect 209 220 214 225
rect 209 218 211 220
rect 213 218 214 220
rect 209 216 214 218
rect 184 212 198 213
rect 184 210 188 212
rect 190 210 198 212
rect 184 209 198 210
rect 169 196 171 198
rect 173 196 181 198
rect 169 192 181 196
rect 193 203 198 209
rect 193 201 194 203
rect 196 201 198 203
rect 193 200 198 201
rect 225 207 230 214
rect 253 229 269 230
rect 253 227 255 229
rect 257 227 269 229
rect 253 225 269 227
rect 265 219 269 225
rect 265 217 266 219
rect 268 217 269 219
rect 280 221 284 230
rect 322 232 327 238
rect 369 236 382 237
rect 369 234 378 236
rect 380 234 382 236
rect 311 229 316 231
rect 280 220 293 221
rect 280 218 285 220
rect 287 218 293 220
rect 280 217 293 218
rect 225 206 227 207
rect 217 205 227 206
rect 229 205 230 207
rect 217 203 230 205
rect 217 201 219 203
rect 221 201 230 203
rect 217 200 230 201
rect 265 197 269 217
rect 287 212 301 213
rect 287 210 295 212
rect 297 210 301 212
rect 287 209 301 210
rect 311 227 312 229
rect 314 227 316 229
rect 311 222 316 227
rect 322 230 324 232
rect 326 230 327 232
rect 369 233 382 234
rect 322 229 327 230
rect 322 228 335 229
rect 322 226 332 228
rect 334 226 335 228
rect 322 225 335 226
rect 311 220 312 222
rect 314 220 316 222
rect 311 218 316 220
rect 287 200 292 209
rect 312 204 316 218
rect 312 202 313 204
rect 315 202 316 204
rect 312 198 316 202
rect 245 196 269 197
rect 245 194 247 196
rect 249 194 269 196
rect 245 193 269 194
rect 304 196 312 198
rect 314 196 316 198
rect 304 192 316 196
rect 336 212 342 214
rect 336 210 337 212
rect 339 210 342 212
rect 336 205 342 210
rect 329 204 342 205
rect 329 202 330 204
rect 332 202 342 204
rect 354 220 366 222
rect 354 218 355 220
rect 357 218 366 220
rect 354 217 366 218
rect 354 216 364 217
rect 362 215 364 216
rect 362 208 366 215
rect 378 212 382 233
rect 378 210 379 212
rect 381 210 382 212
rect 329 201 342 202
rect 378 200 382 210
rect 377 198 382 200
rect 377 196 378 198
rect 380 196 382 198
rect 377 194 382 196
rect 378 192 382 194
rect 389 236 402 237
rect 389 234 391 236
rect 393 234 402 236
rect 389 233 402 234
rect 389 200 393 233
rect 444 232 449 238
rect 444 230 445 232
rect 447 230 449 232
rect 444 229 449 230
rect 436 225 449 229
rect 456 236 469 237
rect 456 234 458 236
rect 460 234 469 236
rect 456 233 469 234
rect 405 217 417 222
rect 407 216 417 217
rect 407 215 409 216
rect 405 212 409 215
rect 405 210 406 212
rect 408 210 409 212
rect 405 208 409 210
rect 429 212 435 214
rect 429 210 432 212
rect 434 210 435 212
rect 429 205 435 210
rect 429 204 442 205
rect 429 202 437 204
rect 439 202 442 204
rect 429 201 442 202
rect 389 198 394 200
rect 389 196 391 198
rect 393 196 394 198
rect 389 194 394 196
rect 389 192 393 194
rect 456 204 460 233
rect 511 232 516 238
rect 511 230 512 232
rect 514 230 516 232
rect 511 229 516 230
rect 503 228 516 229
rect 503 226 504 228
rect 506 226 516 228
rect 503 225 516 226
rect 522 237 526 238
rect 522 233 535 237
rect 522 231 524 233
rect 522 226 526 231
rect 522 224 524 226
rect 472 219 484 222
rect 472 217 480 219
rect 482 217 484 219
rect 474 216 484 217
rect 474 215 476 216
rect 456 202 457 204
rect 459 202 460 204
rect 472 208 476 215
rect 456 200 460 202
rect 496 212 502 214
rect 496 210 499 212
rect 501 210 502 212
rect 496 205 502 210
rect 496 204 509 205
rect 496 202 505 204
rect 507 202 509 204
rect 496 201 509 202
rect 456 198 461 200
rect 456 196 458 198
rect 460 196 461 198
rect 456 194 461 196
rect 456 192 460 194
rect 522 220 526 224
rect 522 218 523 220
rect 525 218 526 220
rect 522 205 526 218
rect 554 221 558 230
rect 537 219 558 221
rect 537 217 551 219
rect 553 217 558 219
rect 564 229 580 230
rect 564 227 576 229
rect 578 227 580 229
rect 564 225 580 227
rect 522 203 527 205
rect 522 201 524 203
rect 526 201 527 203
rect 522 199 527 201
rect 537 212 558 213
rect 537 210 541 212
rect 543 210 558 212
rect 537 209 558 210
rect 554 200 558 209
rect 564 204 568 225
rect 612 232 624 238
rect 564 202 565 204
rect 567 202 568 204
rect 564 197 568 202
rect 603 207 608 214
rect 619 220 624 232
rect 619 218 620 220
rect 622 218 624 220
rect 619 216 624 218
rect 603 205 604 207
rect 606 206 608 207
rect 606 205 616 206
rect 603 200 616 205
rect 564 196 588 197
rect 564 194 584 196
rect 586 194 588 196
rect 564 193 588 194
rect 2 186 632 187
rect 2 184 9 186
rect 11 184 58 186
rect 60 184 68 186
rect 70 184 98 186
rect 100 184 151 186
rect 153 184 172 186
rect 174 184 182 186
rect 184 184 212 186
rect 214 184 265 186
rect 267 184 301 186
rect 303 184 311 186
rect 313 184 525 186
rect 527 184 566 186
rect 568 184 619 186
rect 621 184 632 186
rect 2 174 632 184
rect 2 172 9 174
rect 11 172 58 174
rect 60 172 68 174
rect 70 172 98 174
rect 100 172 151 174
rect 153 172 172 174
rect 174 172 182 174
rect 184 172 212 174
rect 214 172 265 174
rect 267 172 301 174
rect 303 172 311 174
rect 313 172 525 174
rect 527 172 566 174
rect 568 172 619 174
rect 621 172 632 174
rect 2 171 632 172
rect 55 162 67 166
rect 55 160 57 162
rect 59 160 67 162
rect 131 164 155 165
rect 6 157 11 159
rect 6 155 8 157
rect 10 155 11 157
rect 6 153 11 155
rect 6 149 10 153
rect 6 147 7 149
rect 9 147 10 149
rect 6 134 10 147
rect 38 149 42 158
rect 6 132 8 134
rect 6 127 10 132
rect 6 125 8 127
rect 21 148 42 149
rect 21 146 25 148
rect 27 146 39 148
rect 41 146 42 148
rect 21 145 42 146
rect 21 139 35 141
rect 37 139 42 141
rect 21 137 42 139
rect 38 135 42 137
rect 55 140 59 160
rect 131 162 133 164
rect 135 162 155 164
rect 131 161 155 162
rect 79 157 84 158
rect 79 155 80 157
rect 82 155 84 157
rect 79 149 84 155
rect 55 138 60 140
rect 55 136 57 138
rect 59 136 60 138
rect 55 135 60 136
rect 38 131 60 135
rect 38 128 42 131
rect 55 129 57 131
rect 59 129 60 131
rect 70 148 84 149
rect 70 146 74 148
rect 76 146 84 148
rect 70 145 84 146
rect 103 157 116 158
rect 103 155 105 157
rect 107 155 116 157
rect 103 153 116 155
rect 103 152 113 153
rect 111 151 113 152
rect 115 151 116 153
rect 78 140 91 141
rect 78 138 84 140
rect 86 138 91 140
rect 78 137 91 138
rect 55 127 60 129
rect 6 121 19 125
rect 6 120 10 121
rect 87 133 91 137
rect 87 131 88 133
rect 90 131 91 133
rect 87 128 91 131
rect 95 140 100 142
rect 95 138 97 140
rect 99 138 100 140
rect 95 133 100 138
rect 111 144 116 151
rect 151 156 155 161
rect 151 154 152 156
rect 154 154 155 156
rect 95 131 97 133
rect 99 131 100 133
rect 95 126 100 131
rect 95 120 107 126
rect 151 133 155 154
rect 139 131 155 133
rect 139 129 141 131
rect 143 129 155 131
rect 139 128 155 129
rect 169 162 181 166
rect 169 160 171 162
rect 173 160 181 162
rect 245 164 269 165
rect 169 148 173 160
rect 245 162 247 164
rect 249 162 269 164
rect 245 161 269 162
rect 169 146 170 148
rect 172 146 173 148
rect 169 140 173 146
rect 193 157 198 158
rect 193 155 194 157
rect 196 155 198 157
rect 193 149 198 155
rect 169 138 174 140
rect 169 136 171 138
rect 173 136 174 138
rect 169 131 174 136
rect 169 129 171 131
rect 173 129 174 131
rect 184 148 198 149
rect 184 146 188 148
rect 190 146 198 148
rect 184 145 198 146
rect 217 157 230 158
rect 217 155 219 157
rect 221 155 230 157
rect 217 153 230 155
rect 217 152 227 153
rect 225 151 227 152
rect 229 151 230 153
rect 192 140 205 141
rect 192 138 198 140
rect 200 138 205 140
rect 192 137 205 138
rect 169 127 174 129
rect 201 133 205 137
rect 201 131 202 133
rect 204 131 205 133
rect 201 128 205 131
rect 209 140 214 142
rect 209 138 211 140
rect 213 138 214 140
rect 209 133 214 138
rect 225 144 230 151
rect 209 131 211 133
rect 213 131 214 133
rect 209 126 214 131
rect 209 120 221 126
rect 265 141 269 161
rect 287 149 292 158
rect 304 162 316 166
rect 304 160 312 162
rect 314 160 316 162
rect 287 148 301 149
rect 287 146 295 148
rect 297 146 301 148
rect 287 145 301 146
rect 265 139 266 141
rect 268 139 269 141
rect 265 133 269 139
rect 253 131 269 133
rect 253 129 255 131
rect 257 129 269 131
rect 253 128 269 129
rect 280 140 293 141
rect 280 138 285 140
rect 287 138 293 140
rect 280 137 293 138
rect 280 128 284 137
rect 312 156 316 160
rect 312 154 313 156
rect 315 154 316 156
rect 312 140 316 154
rect 311 138 316 140
rect 311 136 312 138
rect 314 136 316 138
rect 378 164 382 166
rect 377 162 382 164
rect 377 160 378 162
rect 380 160 382 162
rect 377 158 382 160
rect 329 156 342 157
rect 329 154 330 156
rect 332 154 342 156
rect 329 153 342 154
rect 336 148 342 153
rect 336 146 337 148
rect 339 146 342 148
rect 336 144 342 146
rect 362 143 366 150
rect 362 142 364 143
rect 354 141 364 142
rect 354 140 366 141
rect 354 138 355 140
rect 357 138 366 140
rect 354 136 366 138
rect 311 131 316 136
rect 311 129 312 131
rect 314 129 316 131
rect 311 127 316 129
rect 322 132 335 133
rect 322 130 332 132
rect 334 130 335 132
rect 322 129 335 130
rect 322 128 327 129
rect 378 148 382 158
rect 378 146 379 148
rect 381 146 382 148
rect 322 126 324 128
rect 326 126 327 128
rect 322 120 327 126
rect 378 125 382 146
rect 369 124 382 125
rect 369 122 378 124
rect 380 122 382 124
rect 369 121 382 122
rect 389 164 393 166
rect 389 162 394 164
rect 389 160 391 162
rect 393 160 394 162
rect 456 164 460 166
rect 389 158 394 160
rect 389 125 393 158
rect 429 156 442 157
rect 405 148 409 150
rect 405 146 406 148
rect 408 146 409 148
rect 405 143 409 146
rect 407 142 409 143
rect 407 141 417 142
rect 405 136 417 141
rect 429 154 437 156
rect 439 154 442 156
rect 429 153 442 154
rect 429 148 435 153
rect 429 146 432 148
rect 434 146 435 148
rect 429 144 435 146
rect 456 162 461 164
rect 456 160 458 162
rect 460 160 461 162
rect 564 164 588 165
rect 456 158 461 160
rect 456 156 460 158
rect 456 154 457 156
rect 459 154 460 156
rect 496 156 509 157
rect 436 129 449 133
rect 444 128 449 129
rect 389 124 402 125
rect 444 126 445 128
rect 447 126 449 128
rect 389 122 391 124
rect 393 122 402 124
rect 389 121 402 122
rect 444 120 449 126
rect 456 125 460 154
rect 472 143 476 150
rect 474 142 476 143
rect 474 141 484 142
rect 472 139 480 141
rect 482 139 484 141
rect 472 136 484 139
rect 496 154 505 156
rect 507 154 509 156
rect 496 153 509 154
rect 496 148 502 153
rect 496 146 499 148
rect 501 146 502 148
rect 496 144 502 146
rect 564 162 584 164
rect 586 162 588 164
rect 564 161 588 162
rect 522 157 527 159
rect 522 155 524 157
rect 526 155 527 157
rect 522 153 527 155
rect 522 140 526 153
rect 522 138 523 140
rect 525 138 526 140
rect 522 134 526 138
rect 554 149 558 158
rect 503 132 516 133
rect 503 130 504 132
rect 506 130 516 132
rect 503 129 516 130
rect 511 128 516 129
rect 456 124 469 125
rect 511 126 512 128
rect 514 126 516 128
rect 456 122 458 124
rect 460 122 469 124
rect 456 121 469 122
rect 511 120 516 126
rect 522 132 524 134
rect 522 127 526 132
rect 522 125 524 127
rect 537 148 558 149
rect 537 146 541 148
rect 543 146 558 148
rect 537 145 558 146
rect 564 156 568 161
rect 564 154 565 156
rect 567 154 568 156
rect 537 139 551 141
rect 553 139 558 141
rect 537 137 558 139
rect 554 128 558 137
rect 564 133 568 154
rect 603 153 616 158
rect 603 151 604 153
rect 606 152 616 153
rect 606 151 608 152
rect 564 131 580 133
rect 564 129 576 131
rect 578 129 580 131
rect 564 128 580 129
rect 603 144 608 151
rect 619 140 624 142
rect 619 138 620 140
rect 622 138 624 140
rect 522 121 535 125
rect 619 126 624 138
rect 522 120 526 121
rect 612 120 624 126
rect 2 114 632 115
rect 2 112 9 114
rect 11 112 58 114
rect 60 112 131 114
rect 133 112 172 114
rect 174 112 245 114
rect 247 112 311 114
rect 313 112 525 114
rect 527 112 586 114
rect 588 112 632 114
rect 2 102 632 112
rect 2 100 9 102
rect 11 100 58 102
rect 60 100 131 102
rect 133 100 172 102
rect 174 100 245 102
rect 247 100 311 102
rect 313 100 525 102
rect 527 100 586 102
rect 588 100 632 102
rect 2 99 632 100
rect 6 93 10 94
rect 6 89 19 93
rect 6 87 8 89
rect 6 82 10 87
rect 6 80 8 82
rect 6 77 10 80
rect 38 83 42 86
rect 55 85 60 87
rect 55 83 57 85
rect 59 83 60 85
rect 95 88 107 94
rect 6 75 7 77
rect 9 75 10 77
rect 6 61 10 75
rect 38 79 60 83
rect 38 77 42 79
rect 21 75 42 77
rect 21 73 35 75
rect 37 73 42 75
rect 55 78 60 79
rect 55 76 57 78
rect 59 76 60 78
rect 55 74 60 76
rect 87 83 91 86
rect 87 81 88 83
rect 90 81 91 83
rect 6 59 11 61
rect 6 57 8 59
rect 10 57 11 59
rect 6 55 11 57
rect 21 68 42 69
rect 21 66 25 68
rect 27 66 39 68
rect 41 66 42 68
rect 21 65 42 66
rect 38 56 42 65
rect 55 54 59 74
rect 87 77 91 81
rect 78 76 91 77
rect 78 74 84 76
rect 86 74 91 76
rect 78 73 91 74
rect 95 83 100 88
rect 95 81 97 83
rect 99 81 100 83
rect 95 76 100 81
rect 95 74 97 76
rect 99 74 100 76
rect 95 72 100 74
rect 70 68 84 69
rect 70 66 74 68
rect 76 66 84 68
rect 70 65 84 66
rect 55 52 57 54
rect 59 52 67 54
rect 55 48 67 52
rect 79 59 84 65
rect 79 57 80 59
rect 82 57 84 59
rect 79 56 84 57
rect 111 63 116 70
rect 139 85 155 86
rect 139 83 141 85
rect 143 83 155 85
rect 139 81 155 83
rect 111 62 113 63
rect 103 61 113 62
rect 115 61 116 63
rect 103 59 116 61
rect 103 57 105 59
rect 107 57 116 59
rect 103 56 116 57
rect 151 60 155 81
rect 151 58 152 60
rect 154 58 155 60
rect 151 53 155 58
rect 131 52 155 53
rect 131 50 133 52
rect 135 50 155 52
rect 131 49 155 50
rect 169 85 174 87
rect 169 83 171 85
rect 173 83 174 85
rect 209 88 221 94
rect 169 78 174 83
rect 169 76 171 78
rect 173 76 174 78
rect 169 74 174 76
rect 201 83 205 86
rect 201 81 202 83
rect 204 81 205 83
rect 169 68 173 74
rect 169 66 170 68
rect 172 66 173 68
rect 169 54 173 66
rect 201 77 205 81
rect 192 76 205 77
rect 192 74 198 76
rect 200 74 205 76
rect 192 73 205 74
rect 209 83 214 88
rect 209 81 211 83
rect 213 81 214 83
rect 209 76 214 81
rect 209 74 211 76
rect 213 74 214 76
rect 209 72 214 74
rect 184 68 198 69
rect 184 66 188 68
rect 190 66 198 68
rect 184 65 198 66
rect 169 52 171 54
rect 173 52 181 54
rect 169 48 181 52
rect 193 59 198 65
rect 193 57 194 59
rect 196 57 198 59
rect 193 56 198 57
rect 225 63 230 70
rect 253 85 269 86
rect 253 83 255 85
rect 257 83 269 85
rect 253 81 269 83
rect 265 75 269 81
rect 265 73 266 75
rect 268 73 269 75
rect 280 77 284 86
rect 322 88 327 94
rect 369 92 382 93
rect 369 90 378 92
rect 380 90 382 92
rect 311 85 316 87
rect 280 76 293 77
rect 280 74 285 76
rect 287 74 293 76
rect 280 73 293 74
rect 225 62 227 63
rect 217 61 227 62
rect 229 61 230 63
rect 217 59 230 61
rect 217 57 219 59
rect 221 57 230 59
rect 217 56 230 57
rect 265 53 269 73
rect 287 68 301 69
rect 287 66 295 68
rect 297 66 301 68
rect 287 65 301 66
rect 311 83 312 85
rect 314 83 316 85
rect 311 78 316 83
rect 322 86 324 88
rect 326 86 327 88
rect 369 89 382 90
rect 322 85 327 86
rect 322 84 335 85
rect 322 82 332 84
rect 334 82 335 84
rect 322 81 335 82
rect 311 76 312 78
rect 314 76 316 78
rect 311 74 316 76
rect 287 56 292 65
rect 312 60 316 74
rect 312 58 313 60
rect 315 58 316 60
rect 312 54 316 58
rect 245 52 269 53
rect 245 50 247 52
rect 249 50 269 52
rect 245 49 269 50
rect 304 52 312 54
rect 314 52 316 54
rect 304 48 316 52
rect 336 68 342 70
rect 336 66 337 68
rect 339 66 342 68
rect 336 61 342 66
rect 329 60 342 61
rect 329 58 330 60
rect 332 58 342 60
rect 354 76 366 78
rect 354 74 355 76
rect 357 74 366 76
rect 354 73 366 74
rect 354 72 364 73
rect 362 71 364 72
rect 362 64 366 71
rect 378 68 382 89
rect 378 66 379 68
rect 381 66 382 68
rect 329 57 342 58
rect 378 56 382 66
rect 377 54 382 56
rect 377 52 378 54
rect 380 52 382 54
rect 377 50 382 52
rect 378 48 382 50
rect 389 92 402 93
rect 389 90 391 92
rect 393 90 402 92
rect 389 89 402 90
rect 389 56 393 89
rect 444 88 449 94
rect 444 86 445 88
rect 447 86 449 88
rect 444 85 449 86
rect 436 81 449 85
rect 456 92 469 93
rect 456 90 458 92
rect 460 90 469 92
rect 456 89 469 90
rect 405 73 417 78
rect 407 72 417 73
rect 407 71 409 72
rect 405 68 409 71
rect 405 66 406 68
rect 408 66 409 68
rect 405 64 409 66
rect 429 68 435 70
rect 429 66 432 68
rect 434 66 435 68
rect 429 61 435 66
rect 429 60 442 61
rect 429 58 437 60
rect 439 58 442 60
rect 429 57 442 58
rect 389 54 394 56
rect 389 52 391 54
rect 393 52 394 54
rect 389 50 394 52
rect 389 48 393 50
rect 456 60 460 89
rect 511 88 516 94
rect 511 86 512 88
rect 514 86 516 88
rect 511 85 516 86
rect 503 84 516 85
rect 503 82 504 84
rect 506 82 516 84
rect 503 81 516 82
rect 522 93 526 94
rect 522 89 535 93
rect 522 87 524 89
rect 522 82 526 87
rect 522 80 524 82
rect 472 75 484 78
rect 472 73 480 75
rect 482 73 484 75
rect 474 72 484 73
rect 474 71 476 72
rect 456 58 457 60
rect 459 58 460 60
rect 472 64 476 71
rect 456 56 460 58
rect 496 68 502 70
rect 496 66 499 68
rect 501 66 502 68
rect 496 61 502 66
rect 496 60 509 61
rect 496 58 505 60
rect 507 58 509 60
rect 496 57 509 58
rect 456 54 461 56
rect 456 52 458 54
rect 460 52 461 54
rect 456 50 461 52
rect 456 48 460 50
rect 522 76 526 80
rect 522 74 523 76
rect 525 74 526 76
rect 522 61 526 74
rect 554 77 558 86
rect 537 75 558 77
rect 537 73 551 75
rect 553 73 558 75
rect 564 85 580 86
rect 564 83 576 85
rect 578 83 580 85
rect 564 81 580 83
rect 522 59 527 61
rect 522 57 524 59
rect 526 57 527 59
rect 522 55 527 57
rect 537 68 558 69
rect 537 66 541 68
rect 543 66 558 68
rect 537 65 558 66
rect 554 56 558 65
rect 564 60 568 81
rect 612 88 624 94
rect 564 58 565 60
rect 567 58 568 60
rect 564 53 568 58
rect 603 63 608 70
rect 619 76 624 88
rect 619 74 620 76
rect 622 74 624 76
rect 619 72 624 74
rect 603 61 604 63
rect 606 62 608 63
rect 606 61 616 62
rect 603 56 616 61
rect 564 52 588 53
rect 564 50 584 52
rect 586 50 588 52
rect 564 49 588 50
rect 2 42 632 43
rect 2 40 9 42
rect 11 40 58 42
rect 60 40 68 42
rect 70 40 98 42
rect 100 40 151 42
rect 153 40 172 42
rect 174 40 182 42
rect 184 40 212 42
rect 214 40 265 42
rect 267 40 301 42
rect 303 40 311 42
rect 313 40 525 42
rect 527 40 566 42
rect 568 40 619 42
rect 621 40 632 42
rect 2 35 632 40
<< alu2 >>
rect 79 301 111 302
rect 79 299 80 301
rect 82 299 105 301
rect 107 299 111 301
rect 79 297 111 299
rect 151 301 225 302
rect 151 300 194 301
rect 151 298 152 300
rect 154 299 194 300
rect 196 299 219 301
rect 221 299 225 301
rect 154 298 225 299
rect 151 297 225 298
rect 312 300 333 301
rect 312 298 313 300
rect 315 298 330 300
rect 332 298 333 300
rect 312 297 333 298
rect 436 300 460 301
rect 436 298 437 300
rect 439 298 457 300
rect 459 298 460 300
rect 436 297 460 298
rect 504 300 568 301
rect 504 298 505 300
rect 507 298 565 300
rect 567 298 568 300
rect 504 297 568 298
rect 38 292 173 293
rect 38 290 39 292
rect 41 290 170 292
rect 172 290 173 292
rect 38 289 173 290
rect 378 292 409 293
rect 378 290 379 292
rect 381 290 406 292
rect 408 290 409 292
rect 378 289 409 290
rect 265 285 359 286
rect 265 283 266 285
rect 268 284 359 285
rect 268 283 355 284
rect 265 282 355 283
rect 357 282 359 284
rect 265 281 359 282
rect 479 285 526 286
rect 479 283 480 285
rect 482 284 526 285
rect 482 283 523 284
rect 479 282 523 283
rect 525 282 526 284
rect 479 281 526 282
rect 87 277 100 278
rect 87 275 88 277
rect 90 275 97 277
rect 99 275 100 277
rect 87 274 100 275
rect 201 277 214 278
rect 201 275 202 277
rect 204 275 211 277
rect 213 275 214 277
rect 201 274 214 275
rect 331 276 508 277
rect 331 274 332 276
rect 334 274 504 276
rect 506 274 508 276
rect 6 247 10 251
rect 201 247 205 274
rect 331 273 508 274
rect 6 243 205 247
rect 6 221 10 243
rect 331 228 508 229
rect 87 227 100 228
rect 87 225 88 227
rect 90 225 97 227
rect 99 225 100 227
rect 87 224 100 225
rect 201 227 214 228
rect 201 225 202 227
rect 204 225 211 227
rect 213 225 214 227
rect 331 226 332 228
rect 334 226 504 228
rect 506 226 508 228
rect 331 225 508 226
rect 201 224 214 225
rect 6 219 7 221
rect 9 219 10 221
rect 6 218 10 219
rect 201 217 205 224
rect 265 220 359 221
rect 265 219 355 220
rect 265 217 266 219
rect 268 218 355 219
rect 357 218 359 220
rect 268 217 359 218
rect 201 213 255 217
rect 265 216 359 217
rect 479 220 526 221
rect 479 219 523 220
rect 479 217 480 219
rect 482 218 523 219
rect 525 218 526 220
rect 482 217 526 218
rect 479 216 526 217
rect 38 212 173 213
rect 38 210 39 212
rect 41 210 170 212
rect 172 210 173 212
rect 38 209 173 210
rect 79 203 111 205
rect 79 201 80 203
rect 82 201 105 203
rect 107 201 111 203
rect 79 200 111 201
rect 151 204 225 205
rect 151 202 152 204
rect 154 203 225 204
rect 154 202 194 203
rect 151 201 194 202
rect 196 201 219 203
rect 221 201 225 203
rect 151 200 225 201
rect 250 185 255 213
rect 378 212 409 213
rect 378 210 379 212
rect 381 210 406 212
rect 408 210 409 212
rect 378 209 409 210
rect 312 204 333 205
rect 312 202 313 204
rect 315 202 330 204
rect 332 202 333 204
rect 312 201 333 202
rect 436 204 460 205
rect 436 202 437 204
rect 439 202 457 204
rect 459 202 460 204
rect 436 201 460 202
rect 504 204 568 205
rect 504 202 505 204
rect 507 202 565 204
rect 567 202 568 204
rect 504 201 568 202
rect 6 181 255 185
rect 6 149 11 181
rect 79 157 111 158
rect 79 155 80 157
rect 82 155 105 157
rect 107 155 111 157
rect 79 153 111 155
rect 151 157 225 158
rect 151 156 194 157
rect 151 154 152 156
rect 154 155 194 156
rect 196 155 219 157
rect 221 155 225 157
rect 154 154 225 155
rect 151 153 225 154
rect 312 156 333 157
rect 312 154 313 156
rect 315 154 330 156
rect 332 154 333 156
rect 312 153 333 154
rect 436 156 460 157
rect 436 154 437 156
rect 439 154 457 156
rect 459 154 460 156
rect 436 153 460 154
rect 504 156 568 157
rect 504 154 505 156
rect 507 154 565 156
rect 567 154 568 156
rect 504 153 568 154
rect 6 147 7 149
rect 9 147 11 149
rect 6 145 11 147
rect 38 148 173 149
rect 38 146 39 148
rect 41 146 170 148
rect 172 146 173 148
rect 38 145 173 146
rect 378 148 409 149
rect 378 146 379 148
rect 381 146 406 148
rect 408 146 409 148
rect 378 145 409 146
rect 265 141 359 142
rect 265 139 266 141
rect 268 140 359 141
rect 268 139 355 140
rect 265 138 355 139
rect 357 138 359 140
rect 265 137 359 138
rect 479 141 526 142
rect 479 139 480 141
rect 482 140 526 141
rect 482 139 523 140
rect 479 138 523 139
rect 525 138 526 140
rect 479 137 526 138
rect 87 133 100 134
rect 87 131 88 133
rect 90 131 97 133
rect 99 131 100 133
rect 87 130 100 131
rect 201 133 214 134
rect 201 131 202 133
rect 204 131 211 133
rect 213 131 214 133
rect 201 130 214 131
rect 331 132 508 133
rect 331 130 332 132
rect 334 130 504 132
rect 506 130 508 132
rect 201 113 205 130
rect 331 129 508 130
rect 6 109 205 113
rect 6 77 10 109
rect 331 84 508 85
rect 87 83 100 84
rect 87 81 88 83
rect 90 81 97 83
rect 99 81 100 83
rect 87 80 100 81
rect 201 83 214 84
rect 201 81 202 83
rect 204 81 211 83
rect 213 81 214 83
rect 331 82 332 84
rect 334 82 504 84
rect 506 82 508 84
rect 331 81 508 82
rect 201 80 214 81
rect 6 75 7 77
rect 9 75 10 77
rect 6 74 10 75
rect 265 76 359 77
rect 265 75 355 76
rect 265 73 266 75
rect 268 74 355 75
rect 357 74 359 76
rect 268 73 359 74
rect 265 72 359 73
rect 479 76 526 77
rect 479 75 523 76
rect 479 73 480 75
rect 482 74 523 75
rect 525 74 526 76
rect 482 73 526 74
rect 479 72 526 73
rect 38 68 173 69
rect 38 66 39 68
rect 41 66 170 68
rect 172 66 173 68
rect 38 65 173 66
rect 378 68 409 69
rect 378 66 379 68
rect 381 66 406 68
rect 408 66 409 68
rect 378 65 409 66
rect 79 59 111 61
rect 79 57 80 59
rect 82 57 105 59
rect 107 57 111 59
rect 79 56 111 57
rect 151 60 225 61
rect 151 58 152 60
rect 154 59 225 60
rect 154 58 194 59
rect 151 57 194 58
rect 196 57 219 59
rect 221 57 225 59
rect 312 60 333 61
rect 312 58 313 60
rect 315 58 330 60
rect 332 58 333 60
rect 312 57 333 58
rect 436 60 460 61
rect 436 58 437 60
rect 439 58 457 60
rect 459 58 460 60
rect 436 57 460 58
rect 504 60 568 61
rect 504 58 505 60
rect 507 58 565 60
rect 567 58 568 60
rect 504 57 568 58
rect 151 56 225 57
<< ptie >>
rect 7 318 13 320
rect 7 316 9 318
rect 11 316 13 318
rect 56 318 62 320
rect 56 316 58 318
rect 60 316 62 318
rect 7 314 13 316
rect 56 314 62 316
rect 96 318 102 320
rect 96 316 98 318
rect 100 316 102 318
rect 96 314 102 316
rect 170 318 176 320
rect 170 316 172 318
rect 174 316 176 318
rect 170 314 176 316
rect 210 318 216 320
rect 210 316 212 318
rect 214 316 216 318
rect 210 314 216 316
rect 309 318 315 320
rect 309 316 311 318
rect 313 316 315 318
rect 309 314 315 316
rect 523 318 529 320
rect 523 316 525 318
rect 527 316 529 318
rect 523 314 529 316
rect 617 318 623 320
rect 617 316 619 318
rect 621 316 623 318
rect 617 314 623 316
rect 7 186 13 188
rect 56 186 62 188
rect 7 184 9 186
rect 11 184 13 186
rect 7 182 13 184
rect 56 184 58 186
rect 60 184 62 186
rect 56 182 62 184
rect 96 186 102 188
rect 96 184 98 186
rect 100 184 102 186
rect 96 182 102 184
rect 170 186 176 188
rect 170 184 172 186
rect 174 184 176 186
rect 170 182 176 184
rect 210 186 216 188
rect 210 184 212 186
rect 214 184 216 186
rect 210 182 216 184
rect 309 186 315 188
rect 309 184 311 186
rect 313 184 315 186
rect 309 182 315 184
rect 523 186 529 188
rect 523 184 525 186
rect 527 184 529 186
rect 523 182 529 184
rect 617 186 623 188
rect 617 184 619 186
rect 621 184 623 186
rect 617 182 623 184
rect 7 174 13 176
rect 7 172 9 174
rect 11 172 13 174
rect 56 174 62 176
rect 56 172 58 174
rect 60 172 62 174
rect 7 170 13 172
rect 56 170 62 172
rect 96 174 102 176
rect 96 172 98 174
rect 100 172 102 174
rect 96 170 102 172
rect 170 174 176 176
rect 170 172 172 174
rect 174 172 176 174
rect 170 170 176 172
rect 210 174 216 176
rect 210 172 212 174
rect 214 172 216 174
rect 210 170 216 172
rect 309 174 315 176
rect 309 172 311 174
rect 313 172 315 174
rect 309 170 315 172
rect 523 174 529 176
rect 523 172 525 174
rect 527 172 529 174
rect 523 170 529 172
rect 617 174 623 176
rect 617 172 619 174
rect 621 172 623 174
rect 617 170 623 172
rect 7 42 13 44
rect 56 42 62 44
rect 7 40 9 42
rect 11 40 13 42
rect 7 38 13 40
rect 56 40 58 42
rect 60 40 62 42
rect 56 38 62 40
rect 96 42 102 44
rect 96 40 98 42
rect 100 40 102 42
rect 96 38 102 40
rect 170 42 176 44
rect 170 40 172 42
rect 174 40 176 42
rect 170 38 176 40
rect 210 42 216 44
rect 210 40 212 42
rect 214 40 216 42
rect 210 38 216 40
rect 309 42 315 44
rect 309 40 311 42
rect 313 40 315 42
rect 309 38 315 40
rect 523 42 529 44
rect 523 40 525 42
rect 527 40 529 42
rect 523 38 529 40
rect 617 42 623 44
rect 617 40 619 42
rect 621 40 623 42
rect 617 38 623 40
<< ntie >>
rect 7 258 13 260
rect 7 256 9 258
rect 11 256 13 258
rect 56 258 62 260
rect 7 254 13 256
rect 56 256 58 258
rect 60 256 62 258
rect 129 258 135 260
rect 56 254 62 256
rect 129 256 131 258
rect 133 256 135 258
rect 170 258 176 260
rect 129 254 135 256
rect 170 256 172 258
rect 174 256 176 258
rect 243 258 249 260
rect 170 254 176 256
rect 243 256 245 258
rect 247 256 249 258
rect 309 258 315 260
rect 243 254 249 256
rect 309 256 311 258
rect 313 256 315 258
rect 523 258 529 260
rect 309 254 315 256
rect 523 256 525 258
rect 527 256 529 258
rect 584 258 590 260
rect 523 254 529 256
rect 584 256 586 258
rect 588 256 590 258
rect 584 254 590 256
rect 7 246 13 248
rect 7 244 9 246
rect 11 244 13 246
rect 56 246 62 248
rect 7 242 13 244
rect 56 244 58 246
rect 60 244 62 246
rect 129 246 135 248
rect 56 242 62 244
rect 129 244 131 246
rect 133 244 135 246
rect 170 246 176 248
rect 129 242 135 244
rect 170 244 172 246
rect 174 244 176 246
rect 243 246 249 248
rect 170 242 176 244
rect 243 244 245 246
rect 247 244 249 246
rect 309 246 315 248
rect 243 242 249 244
rect 309 244 311 246
rect 313 244 315 246
rect 523 246 529 248
rect 309 242 315 244
rect 523 244 525 246
rect 527 244 529 246
rect 584 246 590 248
rect 523 242 529 244
rect 584 244 586 246
rect 588 244 590 246
rect 584 242 590 244
rect 7 114 13 116
rect 7 112 9 114
rect 11 112 13 114
rect 56 114 62 116
rect 7 110 13 112
rect 56 112 58 114
rect 60 112 62 114
rect 129 114 135 116
rect 56 110 62 112
rect 129 112 131 114
rect 133 112 135 114
rect 170 114 176 116
rect 129 110 135 112
rect 170 112 172 114
rect 174 112 176 114
rect 243 114 249 116
rect 170 110 176 112
rect 243 112 245 114
rect 247 112 249 114
rect 309 114 315 116
rect 243 110 249 112
rect 309 112 311 114
rect 313 112 315 114
rect 523 114 529 116
rect 309 110 315 112
rect 523 112 525 114
rect 527 112 529 114
rect 584 114 590 116
rect 523 110 529 112
rect 584 112 586 114
rect 588 112 590 114
rect 584 110 590 112
rect 7 102 13 104
rect 7 100 9 102
rect 11 100 13 102
rect 56 102 62 104
rect 7 98 13 100
rect 56 100 58 102
rect 60 100 62 102
rect 129 102 135 104
rect 56 98 62 100
rect 129 100 131 102
rect 133 100 135 102
rect 170 102 176 104
rect 129 98 135 100
rect 170 100 172 102
rect 174 100 176 102
rect 243 102 249 104
rect 170 98 176 100
rect 243 100 245 102
rect 247 100 249 102
rect 309 102 315 104
rect 243 98 249 100
rect 309 100 311 102
rect 313 100 315 102
rect 523 102 529 104
rect 309 98 315 100
rect 523 100 525 102
rect 527 100 529 102
rect 584 102 590 104
rect 523 98 529 100
rect 584 100 586 102
rect 588 100 590 102
rect 584 98 590 100
<< nmos >>
rect 13 297 15 306
rect 23 297 25 303
rect 33 297 35 303
rect 62 299 64 308
rect 75 299 77 310
rect 82 299 84 310
rect 102 297 104 306
rect 118 302 120 311
rect 128 302 130 311
rect 138 302 140 314
rect 145 302 147 314
rect 176 299 178 308
rect 189 299 191 310
rect 196 299 198 310
rect 216 297 218 306
rect 232 302 234 311
rect 242 302 244 311
rect 252 302 254 314
rect 259 302 261 314
rect 287 299 289 310
rect 294 299 296 310
rect 307 299 309 308
rect 329 303 331 309
rect 339 303 341 311
rect 346 303 348 311
rect 356 303 358 311
rect 363 303 365 311
rect 373 302 375 311
rect 396 302 398 311
rect 406 303 408 311
rect 413 303 415 311
rect 423 303 425 311
rect 430 303 432 311
rect 440 303 442 309
rect 463 302 465 311
rect 473 303 475 311
rect 480 303 482 311
rect 490 303 492 311
rect 497 303 499 311
rect 507 303 509 309
rect 529 297 531 306
rect 539 297 541 303
rect 549 297 551 303
rect 572 302 574 314
rect 579 302 581 314
rect 589 302 591 311
rect 599 302 601 311
rect 615 297 617 306
rect 13 196 15 205
rect 23 199 25 205
rect 33 199 35 205
rect 62 194 64 203
rect 75 192 77 203
rect 82 192 84 203
rect 102 196 104 205
rect 118 191 120 200
rect 128 191 130 200
rect 138 188 140 200
rect 145 188 147 200
rect 176 194 178 203
rect 189 192 191 203
rect 196 192 198 203
rect 216 196 218 205
rect 232 191 234 200
rect 242 191 244 200
rect 252 188 254 200
rect 259 188 261 200
rect 287 192 289 203
rect 294 192 296 203
rect 307 194 309 203
rect 329 193 331 199
rect 339 191 341 199
rect 346 191 348 199
rect 356 191 358 199
rect 363 191 365 199
rect 373 191 375 200
rect 396 191 398 200
rect 406 191 408 199
rect 413 191 415 199
rect 423 191 425 199
rect 430 191 432 199
rect 440 193 442 199
rect 463 191 465 200
rect 473 191 475 199
rect 480 191 482 199
rect 490 191 492 199
rect 497 191 499 199
rect 507 193 509 199
rect 529 196 531 205
rect 539 199 541 205
rect 549 199 551 205
rect 572 188 574 200
rect 579 188 581 200
rect 589 191 591 200
rect 599 191 601 200
rect 615 196 617 205
rect 13 153 15 162
rect 23 153 25 159
rect 33 153 35 159
rect 62 155 64 164
rect 75 155 77 166
rect 82 155 84 166
rect 102 153 104 162
rect 118 158 120 167
rect 128 158 130 167
rect 138 158 140 170
rect 145 158 147 170
rect 176 155 178 164
rect 189 155 191 166
rect 196 155 198 166
rect 216 153 218 162
rect 232 158 234 167
rect 242 158 244 167
rect 252 158 254 170
rect 259 158 261 170
rect 287 155 289 166
rect 294 155 296 166
rect 307 155 309 164
rect 329 159 331 165
rect 339 159 341 167
rect 346 159 348 167
rect 356 159 358 167
rect 363 159 365 167
rect 373 158 375 167
rect 396 158 398 167
rect 406 159 408 167
rect 413 159 415 167
rect 423 159 425 167
rect 430 159 432 167
rect 440 159 442 165
rect 463 158 465 167
rect 473 159 475 167
rect 480 159 482 167
rect 490 159 492 167
rect 497 159 499 167
rect 507 159 509 165
rect 529 153 531 162
rect 539 153 541 159
rect 549 153 551 159
rect 572 158 574 170
rect 579 158 581 170
rect 589 158 591 167
rect 599 158 601 167
rect 615 153 617 162
rect 13 52 15 61
rect 23 55 25 61
rect 33 55 35 61
rect 62 50 64 59
rect 75 48 77 59
rect 82 48 84 59
rect 102 52 104 61
rect 118 47 120 56
rect 128 47 130 56
rect 138 44 140 56
rect 145 44 147 56
rect 176 50 178 59
rect 189 48 191 59
rect 196 48 198 59
rect 216 52 218 61
rect 232 47 234 56
rect 242 47 244 56
rect 252 44 254 56
rect 259 44 261 56
rect 287 48 289 59
rect 294 48 296 59
rect 307 50 309 59
rect 329 49 331 55
rect 339 47 341 55
rect 346 47 348 55
rect 356 47 358 55
rect 363 47 365 55
rect 373 47 375 56
rect 396 47 398 56
rect 406 47 408 55
rect 413 47 415 55
rect 423 47 425 55
rect 430 47 432 55
rect 440 49 442 55
rect 463 47 465 56
rect 473 47 475 55
rect 480 47 482 55
rect 490 47 492 55
rect 497 47 499 55
rect 507 49 509 55
rect 529 52 531 61
rect 539 55 541 61
rect 549 55 551 61
rect 572 44 574 56
rect 579 44 581 56
rect 589 47 591 56
rect 599 47 601 56
rect 615 52 617 61
<< pmos >>
rect 13 267 15 285
rect 26 257 28 278
rect 33 257 35 278
rect 62 266 64 284
rect 72 264 74 277
rect 82 264 84 277
rect 110 257 112 284
rect 126 266 128 284
rect 136 266 138 284
rect 146 257 148 284
rect 176 266 178 284
rect 186 264 188 277
rect 196 264 198 277
rect 224 257 226 284
rect 240 266 242 284
rect 250 266 252 284
rect 260 257 262 284
rect 287 264 289 277
rect 297 264 299 277
rect 307 266 309 284
rect 329 277 331 285
rect 339 257 341 273
rect 346 257 348 273
rect 356 257 358 273
rect 363 257 365 273
rect 373 257 375 275
rect 396 257 398 275
rect 440 277 442 285
rect 406 257 408 273
rect 413 257 415 273
rect 423 257 425 273
rect 430 257 432 273
rect 463 257 465 275
rect 507 277 509 285
rect 473 257 475 273
rect 480 257 482 273
rect 490 257 492 273
rect 497 257 499 273
rect 529 267 531 285
rect 542 257 544 278
rect 549 257 551 278
rect 571 257 573 284
rect 581 266 583 284
rect 591 266 593 284
rect 607 257 609 284
rect 13 217 15 235
rect 26 224 28 245
rect 33 224 35 245
rect 62 218 64 236
rect 72 225 74 238
rect 82 225 84 238
rect 110 218 112 245
rect 126 218 128 236
rect 136 218 138 236
rect 146 218 148 245
rect 176 218 178 236
rect 186 225 188 238
rect 196 225 198 238
rect 224 218 226 245
rect 240 218 242 236
rect 250 218 252 236
rect 260 218 262 245
rect 287 225 289 238
rect 297 225 299 238
rect 307 218 309 236
rect 339 229 341 245
rect 346 229 348 245
rect 356 229 358 245
rect 363 229 365 245
rect 329 217 331 225
rect 373 227 375 245
rect 396 227 398 245
rect 406 229 408 245
rect 413 229 415 245
rect 423 229 425 245
rect 430 229 432 245
rect 463 227 465 245
rect 473 229 475 245
rect 480 229 482 245
rect 490 229 492 245
rect 497 229 499 245
rect 440 217 442 225
rect 507 217 509 225
rect 529 217 531 235
rect 542 224 544 245
rect 549 224 551 245
rect 571 218 573 245
rect 581 218 583 236
rect 591 218 593 236
rect 607 218 609 245
rect 13 123 15 141
rect 26 113 28 134
rect 33 113 35 134
rect 62 122 64 140
rect 72 120 74 133
rect 82 120 84 133
rect 110 113 112 140
rect 126 122 128 140
rect 136 122 138 140
rect 146 113 148 140
rect 176 122 178 140
rect 186 120 188 133
rect 196 120 198 133
rect 224 113 226 140
rect 240 122 242 140
rect 250 122 252 140
rect 260 113 262 140
rect 287 120 289 133
rect 297 120 299 133
rect 307 122 309 140
rect 329 133 331 141
rect 339 113 341 129
rect 346 113 348 129
rect 356 113 358 129
rect 363 113 365 129
rect 373 113 375 131
rect 396 113 398 131
rect 440 133 442 141
rect 406 113 408 129
rect 413 113 415 129
rect 423 113 425 129
rect 430 113 432 129
rect 463 113 465 131
rect 507 133 509 141
rect 473 113 475 129
rect 480 113 482 129
rect 490 113 492 129
rect 497 113 499 129
rect 529 123 531 141
rect 542 113 544 134
rect 549 113 551 134
rect 571 113 573 140
rect 581 122 583 140
rect 591 122 593 140
rect 607 113 609 140
rect 13 73 15 91
rect 26 80 28 101
rect 33 80 35 101
rect 62 74 64 92
rect 72 81 74 94
rect 82 81 84 94
rect 110 74 112 101
rect 126 74 128 92
rect 136 74 138 92
rect 146 74 148 101
rect 176 74 178 92
rect 186 81 188 94
rect 196 81 198 94
rect 224 74 226 101
rect 240 74 242 92
rect 250 74 252 92
rect 260 74 262 101
rect 287 81 289 94
rect 297 81 299 94
rect 307 74 309 92
rect 339 85 341 101
rect 346 85 348 101
rect 356 85 358 101
rect 363 85 365 101
rect 329 73 331 81
rect 373 83 375 101
rect 396 83 398 101
rect 406 85 408 101
rect 413 85 415 101
rect 423 85 425 101
rect 430 85 432 101
rect 463 83 465 101
rect 473 85 475 101
rect 480 85 482 101
rect 490 85 492 101
rect 497 85 499 101
rect 440 73 442 81
rect 507 73 509 81
rect 529 73 531 91
rect 542 80 544 101
rect 549 80 551 101
rect 571 74 573 101
rect 581 74 583 92
rect 591 74 593 92
rect 607 74 609 101
<< polyct0 >>
rect 15 290 17 292
rect 64 290 66 292
rect 134 290 136 292
rect 144 289 146 291
rect 178 290 180 292
rect 248 290 250 292
rect 258 289 260 291
rect 305 290 307 292
rect 354 296 356 298
rect 372 295 374 297
rect 397 295 399 297
rect 347 280 349 282
rect 415 296 417 298
rect 422 280 424 282
rect 464 295 466 297
rect 482 296 484 298
rect 489 280 491 282
rect 531 290 533 292
rect 573 289 575 291
rect 583 290 585 292
rect 15 210 17 212
rect 64 210 66 212
rect 134 210 136 212
rect 144 211 146 213
rect 178 210 180 212
rect 248 210 250 212
rect 258 211 260 213
rect 305 210 307 212
rect 347 220 349 222
rect 354 204 356 206
rect 422 220 424 222
rect 372 205 374 207
rect 397 205 399 207
rect 415 204 417 206
rect 489 220 491 222
rect 464 205 466 207
rect 482 204 484 206
rect 531 210 533 212
rect 573 211 575 213
rect 583 210 585 212
rect 15 146 17 148
rect 64 146 66 148
rect 134 146 136 148
rect 144 145 146 147
rect 178 146 180 148
rect 248 146 250 148
rect 258 145 260 147
rect 305 146 307 148
rect 354 152 356 154
rect 372 151 374 153
rect 397 151 399 153
rect 347 136 349 138
rect 415 152 417 154
rect 422 136 424 138
rect 464 151 466 153
rect 482 152 484 154
rect 489 136 491 138
rect 531 146 533 148
rect 573 145 575 147
rect 583 146 585 148
rect 15 66 17 68
rect 64 66 66 68
rect 134 66 136 68
rect 144 67 146 69
rect 178 66 180 68
rect 248 66 250 68
rect 258 67 260 69
rect 305 66 307 68
rect 347 76 349 78
rect 354 60 356 62
rect 422 76 424 78
rect 372 61 374 63
rect 397 61 399 63
rect 415 60 417 62
rect 489 76 491 78
rect 464 61 466 63
rect 482 60 484 62
rect 531 66 533 68
rect 573 67 575 69
rect 583 66 585 68
<< polyct1 >>
rect 25 290 27 292
rect 74 290 76 292
rect 35 283 37 285
rect 113 295 115 297
rect 84 282 86 284
rect 188 290 190 292
rect 97 282 99 284
rect 227 295 229 297
rect 198 282 200 284
rect 295 290 297 292
rect 211 282 213 284
rect 285 282 287 284
rect 337 290 339 292
rect 364 285 366 287
rect 405 285 407 287
rect 432 290 434 292
rect 324 270 326 272
rect 472 285 474 287
rect 499 290 501 292
rect 445 270 447 272
rect 541 290 543 292
rect 512 270 514 272
rect 604 295 606 297
rect 551 283 553 285
rect 620 282 622 284
rect 35 217 37 219
rect 25 210 27 212
rect 84 218 86 220
rect 97 218 99 220
rect 74 210 76 212
rect 198 218 200 220
rect 211 218 213 220
rect 285 218 287 220
rect 113 205 115 207
rect 188 210 190 212
rect 227 205 229 207
rect 324 230 326 232
rect 295 210 297 212
rect 445 230 447 232
rect 337 210 339 212
rect 364 215 366 217
rect 405 215 407 217
rect 512 230 514 232
rect 432 210 434 212
rect 472 215 474 217
rect 499 210 501 212
rect 551 217 553 219
rect 620 218 622 220
rect 541 210 543 212
rect 604 205 606 207
rect 25 146 27 148
rect 74 146 76 148
rect 35 139 37 141
rect 113 151 115 153
rect 84 138 86 140
rect 188 146 190 148
rect 97 138 99 140
rect 227 151 229 153
rect 198 138 200 140
rect 295 146 297 148
rect 211 138 213 140
rect 285 138 287 140
rect 337 146 339 148
rect 364 141 366 143
rect 405 141 407 143
rect 432 146 434 148
rect 324 126 326 128
rect 472 141 474 143
rect 499 146 501 148
rect 445 126 447 128
rect 541 146 543 148
rect 512 126 514 128
rect 604 151 606 153
rect 551 139 553 141
rect 620 138 622 140
rect 35 73 37 75
rect 25 66 27 68
rect 84 74 86 76
rect 97 74 99 76
rect 74 66 76 68
rect 198 74 200 76
rect 211 74 213 76
rect 285 74 287 76
rect 113 61 115 63
rect 188 66 190 68
rect 227 61 229 63
rect 324 86 326 88
rect 295 66 297 68
rect 445 86 447 88
rect 337 66 339 68
rect 364 71 366 73
rect 405 71 407 73
rect 512 86 514 88
rect 432 66 434 68
rect 472 71 474 73
rect 499 66 501 68
rect 551 73 553 75
rect 620 74 622 76
rect 541 66 543 68
rect 604 61 606 63
<< ndifct0 >>
rect 19 312 21 314
rect 38 312 40 314
rect 28 299 30 301
rect 87 306 89 308
rect 111 307 113 309
rect 97 299 99 301
rect 123 304 125 306
rect 201 306 203 308
rect 225 307 227 309
rect 211 299 213 301
rect 237 304 239 306
rect 282 306 284 308
rect 324 305 326 307
rect 334 305 336 307
rect 351 307 353 309
rect 368 307 370 309
rect 401 307 403 309
rect 418 307 420 309
rect 435 305 437 307
rect 445 305 447 307
rect 468 307 470 309
rect 485 307 487 309
rect 535 312 537 314
rect 502 305 504 307
rect 512 305 514 307
rect 554 312 556 314
rect 544 299 546 301
rect 594 304 596 306
rect 606 307 608 309
rect 620 299 622 301
rect 28 201 30 203
rect 19 188 21 190
rect 97 201 99 203
rect 87 194 89 196
rect 111 193 113 195
rect 38 188 40 190
rect 123 196 125 198
rect 211 201 213 203
rect 201 194 203 196
rect 225 193 227 195
rect 237 196 239 198
rect 282 194 284 196
rect 324 195 326 197
rect 334 195 336 197
rect 351 193 353 195
rect 368 193 370 195
rect 401 193 403 195
rect 418 193 420 195
rect 435 195 437 197
rect 445 195 447 197
rect 468 193 470 195
rect 485 193 487 195
rect 502 195 504 197
rect 512 195 514 197
rect 544 201 546 203
rect 535 188 537 190
rect 554 188 556 190
rect 594 196 596 198
rect 620 201 622 203
rect 606 193 608 195
rect 19 168 21 170
rect 38 168 40 170
rect 28 155 30 157
rect 87 162 89 164
rect 111 163 113 165
rect 97 155 99 157
rect 123 160 125 162
rect 201 162 203 164
rect 225 163 227 165
rect 211 155 213 157
rect 237 160 239 162
rect 282 162 284 164
rect 324 161 326 163
rect 334 161 336 163
rect 351 163 353 165
rect 368 163 370 165
rect 401 163 403 165
rect 418 163 420 165
rect 435 161 437 163
rect 445 161 447 163
rect 468 163 470 165
rect 485 163 487 165
rect 535 168 537 170
rect 502 161 504 163
rect 512 161 514 163
rect 554 168 556 170
rect 544 155 546 157
rect 594 160 596 162
rect 606 163 608 165
rect 620 155 622 157
rect 28 57 30 59
rect 19 44 21 46
rect 97 57 99 59
rect 87 50 89 52
rect 111 49 113 51
rect 38 44 40 46
rect 123 52 125 54
rect 211 57 213 59
rect 201 50 203 52
rect 225 49 227 51
rect 237 52 239 54
rect 282 50 284 52
rect 324 51 326 53
rect 334 51 336 53
rect 351 49 353 51
rect 368 49 370 51
rect 401 49 403 51
rect 418 49 420 51
rect 435 51 437 53
rect 445 51 447 53
rect 468 49 470 51
rect 485 49 487 51
rect 502 51 504 53
rect 512 51 514 53
rect 544 57 546 59
rect 535 44 537 46
rect 554 44 556 46
rect 594 52 596 54
rect 620 57 622 59
rect 606 49 608 51
<< ndifct1 >>
rect 68 316 70 318
rect 8 299 10 301
rect 151 316 153 318
rect 182 316 184 318
rect 57 304 59 306
rect 133 306 135 308
rect 265 316 267 318
rect 301 316 303 318
rect 171 304 173 306
rect 247 306 249 308
rect 312 304 314 306
rect 378 304 380 306
rect 391 304 393 306
rect 458 304 460 306
rect 566 316 568 318
rect 524 299 526 301
rect 584 306 586 308
rect 8 201 10 203
rect 57 196 59 198
rect 133 194 135 196
rect 68 184 70 186
rect 171 196 173 198
rect 151 184 153 186
rect 247 194 249 196
rect 182 184 184 186
rect 312 196 314 198
rect 265 184 267 186
rect 301 184 303 186
rect 378 196 380 198
rect 391 196 393 198
rect 458 196 460 198
rect 524 201 526 203
rect 584 194 586 196
rect 566 184 568 186
rect 68 172 70 174
rect 8 155 10 157
rect 151 172 153 174
rect 182 172 184 174
rect 57 160 59 162
rect 133 162 135 164
rect 265 172 267 174
rect 301 172 303 174
rect 171 160 173 162
rect 247 162 249 164
rect 312 160 314 162
rect 378 160 380 162
rect 391 160 393 162
rect 458 160 460 162
rect 566 172 568 174
rect 524 155 526 157
rect 584 162 586 164
rect 8 57 10 59
rect 57 52 59 54
rect 133 50 135 52
rect 68 40 70 42
rect 171 52 173 54
rect 151 40 153 42
rect 247 50 249 52
rect 182 40 184 42
rect 312 52 314 54
rect 265 40 267 42
rect 301 40 303 42
rect 378 52 380 54
rect 391 52 393 54
rect 458 52 460 54
rect 524 57 526 59
rect 584 50 586 52
rect 566 40 568 42
<< ntiect1 >>
rect 9 256 11 258
rect 58 256 60 258
rect 131 256 133 258
rect 172 256 174 258
rect 245 256 247 258
rect 311 256 313 258
rect 525 256 527 258
rect 586 256 588 258
rect 9 244 11 246
rect 58 244 60 246
rect 131 244 133 246
rect 172 244 174 246
rect 245 244 247 246
rect 311 244 313 246
rect 525 244 527 246
rect 586 244 588 246
rect 9 112 11 114
rect 58 112 60 114
rect 131 112 133 114
rect 172 112 174 114
rect 245 112 247 114
rect 311 112 313 114
rect 525 112 527 114
rect 586 112 588 114
rect 9 100 11 102
rect 58 100 60 102
rect 131 100 133 102
rect 172 100 174 102
rect 245 100 247 102
rect 311 100 313 102
rect 525 100 527 102
rect 586 100 588 102
<< ptiect1 >>
rect 9 316 11 318
rect 58 316 60 318
rect 98 316 100 318
rect 172 316 174 318
rect 212 316 214 318
rect 311 316 313 318
rect 525 316 527 318
rect 619 316 621 318
rect 9 184 11 186
rect 58 184 60 186
rect 98 184 100 186
rect 172 184 174 186
rect 212 184 214 186
rect 311 184 313 186
rect 525 184 527 186
rect 619 184 621 186
rect 9 172 11 174
rect 58 172 60 174
rect 98 172 100 174
rect 172 172 174 174
rect 212 172 214 174
rect 311 172 313 174
rect 525 172 527 174
rect 619 172 621 174
rect 9 40 11 42
rect 58 40 60 42
rect 98 40 100 42
rect 172 40 174 42
rect 212 40 214 42
rect 311 40 313 42
rect 525 40 527 42
rect 619 40 621 42
<< pdifct0 >>
rect 19 259 21 261
rect 38 266 40 268
rect 105 280 107 282
rect 67 268 69 270
rect 77 273 79 275
rect 77 266 79 268
rect 87 266 89 268
rect 115 266 117 268
rect 131 280 133 282
rect 131 273 133 275
rect 115 259 117 261
rect 151 265 153 267
rect 219 280 221 282
rect 181 268 183 270
rect 191 273 193 275
rect 191 266 193 268
rect 201 266 203 268
rect 229 266 231 268
rect 245 280 247 282
rect 245 273 247 275
rect 229 259 231 261
rect 265 265 267 267
rect 282 266 284 268
rect 292 273 294 275
rect 292 266 294 268
rect 302 268 304 270
rect 324 281 326 283
rect 334 259 336 261
rect 351 269 353 271
rect 368 259 370 261
rect 445 281 447 283
rect 401 259 403 261
rect 418 269 420 271
rect 435 259 437 261
rect 512 281 514 283
rect 468 259 470 261
rect 485 269 487 271
rect 502 259 504 261
rect 535 259 537 261
rect 554 266 556 268
rect 566 265 568 267
rect 586 280 588 282
rect 586 273 588 275
rect 602 266 604 268
rect 602 259 604 261
rect 612 280 614 282
rect 19 241 21 243
rect 38 234 40 236
rect 67 232 69 234
rect 77 234 79 236
rect 77 227 79 229
rect 87 234 89 236
rect 105 220 107 222
rect 115 241 117 243
rect 115 234 117 236
rect 131 227 133 229
rect 131 220 133 222
rect 151 235 153 237
rect 181 232 183 234
rect 191 234 193 236
rect 191 227 193 229
rect 201 234 203 236
rect 219 220 221 222
rect 229 241 231 243
rect 229 234 231 236
rect 245 227 247 229
rect 245 220 247 222
rect 334 241 336 243
rect 265 235 267 237
rect 282 234 284 236
rect 292 234 294 236
rect 292 227 294 229
rect 302 232 304 234
rect 351 231 353 233
rect 368 241 370 243
rect 324 219 326 221
rect 401 241 403 243
rect 418 231 420 233
rect 435 241 437 243
rect 468 241 470 243
rect 485 231 487 233
rect 502 241 504 243
rect 535 241 537 243
rect 445 219 447 221
rect 512 219 514 221
rect 554 234 556 236
rect 566 235 568 237
rect 602 241 604 243
rect 586 227 588 229
rect 586 220 588 222
rect 602 234 604 236
rect 612 220 614 222
rect 19 115 21 117
rect 38 122 40 124
rect 105 136 107 138
rect 67 124 69 126
rect 77 129 79 131
rect 77 122 79 124
rect 87 122 89 124
rect 115 122 117 124
rect 131 136 133 138
rect 131 129 133 131
rect 115 115 117 117
rect 151 121 153 123
rect 219 136 221 138
rect 181 124 183 126
rect 191 129 193 131
rect 191 122 193 124
rect 201 122 203 124
rect 229 122 231 124
rect 245 136 247 138
rect 245 129 247 131
rect 229 115 231 117
rect 265 121 267 123
rect 282 122 284 124
rect 292 129 294 131
rect 292 122 294 124
rect 302 124 304 126
rect 324 137 326 139
rect 334 115 336 117
rect 351 125 353 127
rect 368 115 370 117
rect 445 137 447 139
rect 401 115 403 117
rect 418 125 420 127
rect 435 115 437 117
rect 512 137 514 139
rect 468 115 470 117
rect 485 125 487 127
rect 502 115 504 117
rect 535 115 537 117
rect 554 122 556 124
rect 566 121 568 123
rect 586 136 588 138
rect 586 129 588 131
rect 602 122 604 124
rect 602 115 604 117
rect 612 136 614 138
rect 19 97 21 99
rect 38 90 40 92
rect 67 88 69 90
rect 77 90 79 92
rect 77 83 79 85
rect 87 90 89 92
rect 105 76 107 78
rect 115 97 117 99
rect 115 90 117 92
rect 131 83 133 85
rect 131 76 133 78
rect 151 91 153 93
rect 181 88 183 90
rect 191 90 193 92
rect 191 83 193 85
rect 201 90 203 92
rect 219 76 221 78
rect 229 97 231 99
rect 229 90 231 92
rect 245 83 247 85
rect 245 76 247 78
rect 334 97 336 99
rect 265 91 267 93
rect 282 90 284 92
rect 292 90 294 92
rect 292 83 294 85
rect 302 88 304 90
rect 351 87 353 89
rect 368 97 370 99
rect 324 75 326 77
rect 401 97 403 99
rect 418 87 420 89
rect 435 97 437 99
rect 468 97 470 99
rect 485 87 487 89
rect 502 97 504 99
rect 535 97 537 99
rect 445 75 447 77
rect 512 75 514 77
rect 554 90 556 92
rect 566 91 568 93
rect 602 97 604 99
rect 586 83 588 85
rect 586 76 588 78
rect 602 90 604 92
rect 612 76 614 78
<< pdifct1 >>
rect 8 276 10 278
rect 8 269 10 271
rect 57 280 59 282
rect 57 273 59 275
rect 141 273 143 275
rect 171 280 173 282
rect 171 273 173 275
rect 255 273 257 275
rect 312 280 314 282
rect 312 273 314 275
rect 378 266 380 268
rect 391 266 393 268
rect 458 266 460 268
rect 524 276 526 278
rect 524 269 526 271
rect 576 273 578 275
rect 8 231 10 233
rect 8 224 10 226
rect 57 227 59 229
rect 57 220 59 222
rect 141 227 143 229
rect 171 227 173 229
rect 171 220 173 222
rect 255 227 257 229
rect 312 227 314 229
rect 312 220 314 222
rect 378 234 380 236
rect 391 234 393 236
rect 458 234 460 236
rect 524 231 526 233
rect 524 224 526 226
rect 576 227 578 229
rect 8 132 10 134
rect 8 125 10 127
rect 57 136 59 138
rect 57 129 59 131
rect 141 129 143 131
rect 171 136 173 138
rect 171 129 173 131
rect 255 129 257 131
rect 312 136 314 138
rect 312 129 314 131
rect 378 122 380 124
rect 391 122 393 124
rect 458 122 460 124
rect 524 132 526 134
rect 524 125 526 127
rect 576 129 578 131
rect 8 87 10 89
rect 8 80 10 82
rect 57 83 59 85
rect 57 76 59 78
rect 141 83 143 85
rect 171 83 173 85
rect 171 76 173 78
rect 255 83 257 85
rect 312 83 314 85
rect 312 76 314 78
rect 378 90 380 92
rect 391 90 393 92
rect 458 90 460 92
rect 524 87 526 89
rect 524 80 526 82
rect 576 83 578 85
<< alu0 >>
rect 17 314 23 315
rect 17 312 19 314
rect 21 312 23 314
rect 17 311 23 312
rect 36 314 42 315
rect 36 312 38 314
rect 40 312 42 314
rect 36 311 42 312
rect 109 309 115 315
rect 71 308 91 309
rect 71 306 87 308
rect 89 306 91 308
rect 109 307 111 309
rect 113 307 115 309
rect 109 306 115 307
rect 122 306 126 308
rect 71 305 91 306
rect 14 301 32 302
rect 14 299 28 301
rect 30 299 32 301
rect 14 298 32 299
rect 14 292 18 298
rect 14 290 15 292
rect 17 290 18 292
rect 10 269 11 280
rect 14 277 18 290
rect 33 285 39 286
rect 59 302 60 304
rect 71 301 75 305
rect 122 304 123 306
rect 125 304 126 306
rect 63 297 75 301
rect 63 292 67 297
rect 63 290 64 292
rect 66 290 67 292
rect 14 273 29 277
rect 25 269 29 273
rect 63 278 67 290
rect 96 301 100 303
rect 96 299 97 301
rect 99 299 100 301
rect 96 293 100 299
rect 122 301 126 304
rect 122 297 146 301
rect 96 289 107 293
rect 63 275 80 278
rect 63 274 77 275
rect 76 273 77 274
rect 79 273 80 275
rect 65 270 71 271
rect 25 268 42 269
rect 25 266 38 268
rect 40 266 42 268
rect 25 265 42 266
rect 65 268 67 270
rect 69 268 71 270
rect 17 261 23 262
rect 17 259 19 261
rect 21 259 23 261
rect 65 259 71 268
rect 76 268 80 273
rect 103 283 107 289
rect 142 293 146 297
rect 122 292 138 293
rect 122 290 134 292
rect 136 290 138 292
rect 122 289 138 290
rect 142 291 147 293
rect 142 289 144 291
rect 146 289 147 291
rect 122 283 126 289
rect 142 287 147 289
rect 142 285 146 287
rect 103 282 126 283
rect 103 280 105 282
rect 107 280 126 282
rect 103 279 126 280
rect 76 266 77 268
rect 79 266 80 268
rect 76 264 80 266
rect 85 268 91 269
rect 85 266 87 268
rect 89 266 91 268
rect 85 259 91 266
rect 114 268 118 270
rect 114 266 115 268
rect 117 266 118 268
rect 114 261 118 266
rect 122 268 126 279
rect 130 282 146 285
rect 130 280 131 282
rect 133 281 146 282
rect 133 280 134 281
rect 130 275 134 280
rect 130 273 131 275
rect 133 273 134 275
rect 130 271 134 273
rect 223 309 229 315
rect 185 308 205 309
rect 185 306 201 308
rect 203 306 205 308
rect 223 307 225 309
rect 227 307 229 309
rect 223 306 229 307
rect 236 306 240 308
rect 185 305 205 306
rect 173 302 174 304
rect 185 301 189 305
rect 236 304 237 306
rect 239 304 240 306
rect 280 308 300 309
rect 280 306 282 308
rect 284 306 300 308
rect 280 305 300 306
rect 177 297 189 301
rect 177 292 181 297
rect 177 290 178 292
rect 180 290 181 292
rect 177 278 181 290
rect 210 301 214 303
rect 210 299 211 301
rect 213 299 214 301
rect 210 293 214 299
rect 236 301 240 304
rect 236 297 260 301
rect 210 289 221 293
rect 177 275 194 278
rect 177 274 191 275
rect 190 273 191 274
rect 193 273 194 275
rect 179 270 185 271
rect 179 268 181 270
rect 183 268 185 270
rect 122 267 155 268
rect 122 265 151 267
rect 153 265 155 267
rect 122 264 155 265
rect 114 259 115 261
rect 117 259 118 261
rect 179 259 185 268
rect 190 268 194 273
rect 217 283 221 289
rect 256 293 260 297
rect 236 292 252 293
rect 236 290 248 292
rect 250 290 252 292
rect 236 289 252 290
rect 256 291 261 293
rect 256 289 258 291
rect 260 289 261 291
rect 236 283 240 289
rect 256 287 261 289
rect 256 285 260 287
rect 217 282 240 283
rect 217 280 219 282
rect 221 280 240 282
rect 217 279 240 280
rect 190 266 191 268
rect 193 266 194 268
rect 190 264 194 266
rect 199 268 205 269
rect 199 266 201 268
rect 203 266 205 268
rect 199 259 205 266
rect 228 268 232 270
rect 228 266 229 268
rect 231 266 232 268
rect 228 261 232 266
rect 236 268 240 279
rect 244 282 260 285
rect 244 280 245 282
rect 247 281 260 282
rect 296 301 300 305
rect 311 302 312 304
rect 296 297 308 301
rect 304 292 308 297
rect 304 290 305 292
rect 307 290 308 292
rect 247 280 248 281
rect 244 275 248 280
rect 244 273 245 275
rect 247 273 248 275
rect 244 271 248 273
rect 304 278 308 290
rect 291 275 308 278
rect 291 273 292 275
rect 294 274 308 275
rect 322 307 328 308
rect 322 305 324 307
rect 326 305 328 307
rect 322 304 328 305
rect 332 307 338 315
rect 332 305 334 307
rect 336 305 338 307
rect 349 309 364 310
rect 349 307 351 309
rect 353 307 364 309
rect 349 306 364 307
rect 332 304 338 305
rect 322 284 326 304
rect 360 301 364 306
rect 367 309 371 315
rect 367 307 368 309
rect 370 307 371 309
rect 367 305 371 307
rect 346 298 357 300
rect 346 296 354 298
rect 356 296 357 298
rect 360 299 374 301
rect 360 297 375 299
rect 346 294 357 296
rect 370 295 372 297
rect 374 295 375 297
rect 346 284 350 294
rect 370 293 375 295
rect 322 283 350 284
rect 322 281 324 283
rect 326 282 350 283
rect 326 281 347 282
rect 322 280 347 281
rect 349 280 350 282
rect 366 283 367 289
rect 346 278 350 280
rect 294 273 295 274
rect 280 268 286 269
rect 236 267 269 268
rect 236 265 265 267
rect 267 265 269 267
rect 236 264 269 265
rect 280 266 282 268
rect 284 266 286 268
rect 228 259 229 261
rect 231 259 232 261
rect 280 259 286 266
rect 291 268 295 273
rect 370 276 374 293
rect 358 272 374 276
rect 291 266 292 268
rect 294 266 295 268
rect 291 264 295 266
rect 300 270 306 271
rect 300 268 302 270
rect 304 268 306 270
rect 300 259 306 268
rect 349 271 362 272
rect 349 269 351 271
rect 353 269 362 271
rect 349 268 362 269
rect 400 309 404 315
rect 400 307 401 309
rect 403 307 404 309
rect 400 305 404 307
rect 407 309 422 310
rect 407 307 418 309
rect 420 307 422 309
rect 407 306 422 307
rect 433 307 439 315
rect 467 309 471 315
rect 407 301 411 306
rect 433 305 435 307
rect 437 305 439 307
rect 433 304 439 305
rect 443 307 449 308
rect 443 305 445 307
rect 447 305 449 307
rect 443 304 449 305
rect 397 299 411 301
rect 396 297 411 299
rect 414 298 425 300
rect 396 295 397 297
rect 399 295 401 297
rect 396 293 401 295
rect 414 296 415 298
rect 417 296 425 298
rect 414 294 425 296
rect 397 276 401 293
rect 404 283 405 289
rect 421 284 425 294
rect 445 284 449 304
rect 421 283 449 284
rect 421 282 445 283
rect 421 280 422 282
rect 424 281 445 282
rect 447 281 449 283
rect 424 280 449 281
rect 467 307 468 309
rect 470 307 471 309
rect 467 305 471 307
rect 474 309 489 310
rect 474 307 485 309
rect 487 307 489 309
rect 474 306 489 307
rect 500 307 506 315
rect 533 314 539 315
rect 533 312 535 314
rect 537 312 539 314
rect 533 311 539 312
rect 552 314 558 315
rect 552 312 554 314
rect 556 312 558 314
rect 552 311 558 312
rect 604 309 610 315
rect 474 301 478 306
rect 500 305 502 307
rect 504 305 506 307
rect 500 304 506 305
rect 510 307 516 308
rect 510 305 512 307
rect 514 305 516 307
rect 510 304 516 305
rect 464 299 478 301
rect 421 278 425 280
rect 397 272 413 276
rect 409 271 422 272
rect 409 269 418 271
rect 420 269 422 271
rect 409 268 422 269
rect 463 297 478 299
rect 481 298 492 300
rect 463 295 464 297
rect 466 295 468 297
rect 463 293 468 295
rect 481 296 482 298
rect 484 296 492 298
rect 481 294 492 296
rect 464 276 468 293
rect 471 283 472 289
rect 488 284 492 294
rect 512 284 516 304
rect 593 306 597 308
rect 604 307 606 309
rect 608 307 610 309
rect 604 306 610 307
rect 488 283 516 284
rect 488 282 512 283
rect 488 280 489 282
rect 491 281 512 282
rect 514 281 516 283
rect 491 280 516 281
rect 530 301 548 302
rect 530 299 544 301
rect 546 299 548 301
rect 530 298 548 299
rect 488 278 492 280
rect 530 292 534 298
rect 530 290 531 292
rect 533 290 534 292
rect 464 272 480 276
rect 476 271 489 272
rect 476 269 485 271
rect 487 269 489 271
rect 476 268 489 269
rect 526 269 527 280
rect 530 277 534 290
rect 593 304 594 306
rect 596 304 597 306
rect 593 301 597 304
rect 549 285 555 286
rect 530 273 545 277
rect 541 269 545 273
rect 573 297 597 301
rect 573 293 577 297
rect 619 301 623 303
rect 619 299 620 301
rect 622 299 623 301
rect 572 291 577 293
rect 572 289 573 291
rect 575 289 577 291
rect 581 292 597 293
rect 581 290 583 292
rect 585 290 597 292
rect 581 289 597 290
rect 572 287 577 289
rect 573 285 577 287
rect 573 282 589 285
rect 573 281 586 282
rect 585 280 586 281
rect 588 280 589 282
rect 585 275 589 280
rect 585 273 586 275
rect 588 273 589 275
rect 585 271 589 273
rect 593 283 597 289
rect 619 293 623 299
rect 612 289 623 293
rect 612 283 616 289
rect 593 282 616 283
rect 593 280 612 282
rect 614 280 616 282
rect 593 279 616 280
rect 541 268 558 269
rect 593 268 597 279
rect 541 266 554 268
rect 556 266 558 268
rect 541 265 558 266
rect 564 267 597 268
rect 564 265 566 267
rect 568 265 597 267
rect 564 264 597 265
rect 601 268 605 270
rect 601 266 602 268
rect 604 266 605 268
rect 333 261 337 263
rect 333 259 334 261
rect 336 259 337 261
rect 366 261 372 262
rect 366 259 368 261
rect 370 259 372 261
rect 399 261 405 262
rect 399 259 401 261
rect 403 259 405 261
rect 434 261 438 263
rect 434 259 435 261
rect 437 259 438 261
rect 466 261 472 262
rect 466 259 468 261
rect 470 259 472 261
rect 501 261 505 263
rect 501 259 502 261
rect 504 259 505 261
rect 533 261 539 262
rect 533 259 535 261
rect 537 259 539 261
rect 601 261 605 266
rect 601 259 602 261
rect 604 259 605 261
rect 17 241 19 243
rect 21 241 23 243
rect 17 240 23 241
rect 25 236 42 237
rect 25 234 38 236
rect 40 234 42 236
rect 25 233 42 234
rect 65 234 71 243
rect 10 222 11 233
rect 25 229 29 233
rect 65 232 67 234
rect 69 232 71 234
rect 65 231 71 232
rect 76 236 80 238
rect 76 234 77 236
rect 79 234 80 236
rect 14 225 29 229
rect 76 229 80 234
rect 85 236 91 243
rect 114 241 115 243
rect 117 241 118 243
rect 85 234 87 236
rect 89 234 91 236
rect 85 233 91 234
rect 114 236 118 241
rect 114 234 115 236
rect 117 234 118 236
rect 114 232 118 234
rect 122 237 155 238
rect 122 235 151 237
rect 153 235 155 237
rect 122 234 155 235
rect 179 234 185 243
rect 76 228 77 229
rect 14 212 18 225
rect 63 227 77 228
rect 79 227 80 229
rect 63 224 80 227
rect 33 216 39 217
rect 14 210 15 212
rect 17 210 18 212
rect 14 204 18 210
rect 14 203 32 204
rect 14 201 28 203
rect 30 201 32 203
rect 14 200 32 201
rect 63 212 67 224
rect 122 223 126 234
rect 179 232 181 234
rect 183 232 185 234
rect 179 231 185 232
rect 190 236 194 238
rect 190 234 191 236
rect 193 234 194 236
rect 103 222 126 223
rect 103 220 105 222
rect 107 220 126 222
rect 103 219 126 220
rect 103 213 107 219
rect 63 210 64 212
rect 66 210 67 212
rect 63 205 67 210
rect 63 201 75 205
rect 59 198 60 200
rect 71 197 75 201
rect 96 209 107 213
rect 96 203 100 209
rect 122 213 126 219
rect 130 229 134 231
rect 130 227 131 229
rect 133 227 134 229
rect 130 222 134 227
rect 130 220 131 222
rect 133 221 134 222
rect 133 220 146 221
rect 130 217 146 220
rect 142 215 146 217
rect 142 213 147 215
rect 122 212 138 213
rect 122 210 134 212
rect 136 210 138 212
rect 122 209 138 210
rect 142 211 144 213
rect 146 211 147 213
rect 142 209 147 211
rect 96 201 97 203
rect 99 201 100 203
rect 96 199 100 201
rect 142 205 146 209
rect 122 201 146 205
rect 122 198 126 201
rect 71 196 91 197
rect 122 196 123 198
rect 125 196 126 198
rect 71 194 87 196
rect 89 194 91 196
rect 71 193 91 194
rect 109 195 115 196
rect 109 193 111 195
rect 113 193 115 195
rect 122 194 126 196
rect 190 229 194 234
rect 199 236 205 243
rect 228 241 229 243
rect 231 241 232 243
rect 199 234 201 236
rect 203 234 205 236
rect 199 233 205 234
rect 228 236 232 241
rect 228 234 229 236
rect 231 234 232 236
rect 228 232 232 234
rect 236 237 269 238
rect 236 235 265 237
rect 267 235 269 237
rect 236 234 269 235
rect 280 236 286 243
rect 280 234 282 236
rect 284 234 286 236
rect 190 228 191 229
rect 177 227 191 228
rect 193 227 194 229
rect 177 224 194 227
rect 177 212 181 224
rect 236 223 240 234
rect 280 233 286 234
rect 291 236 295 238
rect 291 234 292 236
rect 294 234 295 236
rect 217 222 240 223
rect 217 220 219 222
rect 221 220 240 222
rect 217 219 240 220
rect 217 213 221 219
rect 177 210 178 212
rect 180 210 181 212
rect 177 205 181 210
rect 177 201 189 205
rect 173 198 174 200
rect 17 190 23 191
rect 17 188 19 190
rect 21 188 23 190
rect 17 187 23 188
rect 36 190 42 191
rect 36 188 38 190
rect 40 188 42 190
rect 36 187 42 188
rect 109 187 115 193
rect 185 197 189 201
rect 210 209 221 213
rect 210 203 214 209
rect 236 213 240 219
rect 244 229 248 231
rect 244 227 245 229
rect 247 227 248 229
rect 244 222 248 227
rect 244 220 245 222
rect 247 221 248 222
rect 247 220 260 221
rect 244 217 260 220
rect 256 215 260 217
rect 291 229 295 234
rect 300 234 306 243
rect 333 241 334 243
rect 336 241 337 243
rect 333 239 337 241
rect 366 241 368 243
rect 370 241 372 243
rect 366 240 372 241
rect 399 241 401 243
rect 403 241 405 243
rect 399 240 405 241
rect 434 241 435 243
rect 437 241 438 243
rect 434 239 438 241
rect 466 241 468 243
rect 470 241 472 243
rect 466 240 472 241
rect 501 241 502 243
rect 504 241 505 243
rect 501 239 505 241
rect 533 241 535 243
rect 537 241 539 243
rect 533 240 539 241
rect 601 241 602 243
rect 604 241 605 243
rect 300 232 302 234
rect 304 232 306 234
rect 300 231 306 232
rect 291 227 292 229
rect 294 228 295 229
rect 294 227 308 228
rect 291 224 308 227
rect 256 213 261 215
rect 236 212 252 213
rect 236 210 248 212
rect 250 210 252 212
rect 236 209 252 210
rect 256 211 258 213
rect 260 211 261 213
rect 256 209 261 211
rect 210 201 211 203
rect 213 201 214 203
rect 210 199 214 201
rect 256 205 260 209
rect 236 201 260 205
rect 236 198 240 201
rect 185 196 205 197
rect 236 196 237 198
rect 239 196 240 198
rect 304 212 308 224
rect 349 233 362 234
rect 349 231 351 233
rect 353 231 362 233
rect 349 230 362 231
rect 358 226 374 230
rect 346 222 350 224
rect 304 210 305 212
rect 307 210 308 212
rect 304 205 308 210
rect 296 201 308 205
rect 296 197 300 201
rect 311 198 312 200
rect 185 194 201 196
rect 203 194 205 196
rect 185 193 205 194
rect 223 195 229 196
rect 223 193 225 195
rect 227 193 229 195
rect 236 194 240 196
rect 280 196 300 197
rect 280 194 282 196
rect 284 194 300 196
rect 280 193 300 194
rect 223 187 229 193
rect 322 221 347 222
rect 322 219 324 221
rect 326 220 347 221
rect 349 220 350 222
rect 326 219 350 220
rect 322 218 350 219
rect 322 198 326 218
rect 346 208 350 218
rect 366 213 367 219
rect 370 209 374 226
rect 346 206 357 208
rect 346 204 354 206
rect 356 204 357 206
rect 370 207 375 209
rect 370 205 372 207
rect 374 205 375 207
rect 346 202 357 204
rect 360 203 375 205
rect 360 201 374 203
rect 322 197 328 198
rect 322 195 324 197
rect 326 195 328 197
rect 322 194 328 195
rect 332 197 338 198
rect 332 195 334 197
rect 336 195 338 197
rect 360 196 364 201
rect 332 187 338 195
rect 349 195 364 196
rect 349 193 351 195
rect 353 193 364 195
rect 349 192 364 193
rect 367 195 371 197
rect 367 193 368 195
rect 370 193 371 195
rect 367 187 371 193
rect 409 233 422 234
rect 409 231 418 233
rect 420 231 422 233
rect 409 230 422 231
rect 397 226 413 230
rect 397 209 401 226
rect 476 233 489 234
rect 421 222 425 224
rect 404 213 405 219
rect 421 220 422 222
rect 424 221 449 222
rect 424 220 445 221
rect 421 219 445 220
rect 447 219 449 221
rect 421 218 449 219
rect 396 207 401 209
rect 421 208 425 218
rect 396 205 397 207
rect 399 205 401 207
rect 414 206 425 208
rect 396 203 411 205
rect 397 201 411 203
rect 414 204 415 206
rect 417 204 425 206
rect 414 202 425 204
rect 400 195 404 197
rect 400 193 401 195
rect 403 193 404 195
rect 400 187 404 193
rect 407 196 411 201
rect 445 198 449 218
rect 433 197 439 198
rect 407 195 422 196
rect 407 193 418 195
rect 420 193 422 195
rect 407 192 422 193
rect 433 195 435 197
rect 437 195 439 197
rect 433 187 439 195
rect 443 197 449 198
rect 443 195 445 197
rect 447 195 449 197
rect 443 194 449 195
rect 476 231 485 233
rect 487 231 489 233
rect 476 230 489 231
rect 464 226 480 230
rect 464 209 468 226
rect 564 237 597 238
rect 541 236 558 237
rect 541 234 554 236
rect 556 234 558 236
rect 564 235 566 237
rect 568 235 597 237
rect 564 234 597 235
rect 541 233 558 234
rect 488 222 492 224
rect 471 213 472 219
rect 488 220 489 222
rect 491 221 516 222
rect 491 220 512 221
rect 488 219 512 220
rect 514 219 516 221
rect 488 218 516 219
rect 463 207 468 209
rect 488 208 492 218
rect 463 205 464 207
rect 466 205 468 207
rect 481 206 492 208
rect 463 203 478 205
rect 464 201 478 203
rect 481 204 482 206
rect 484 204 492 206
rect 481 202 492 204
rect 467 195 471 197
rect 467 193 468 195
rect 470 193 471 195
rect 467 187 471 193
rect 474 196 478 201
rect 512 198 516 218
rect 526 222 527 233
rect 541 229 545 233
rect 530 225 545 229
rect 530 212 534 225
rect 585 229 589 231
rect 585 227 586 229
rect 588 227 589 229
rect 549 216 555 217
rect 530 210 531 212
rect 533 210 534 212
rect 530 204 534 210
rect 530 203 548 204
rect 530 201 544 203
rect 546 201 548 203
rect 530 200 548 201
rect 585 222 589 227
rect 585 221 586 222
rect 573 220 586 221
rect 588 220 589 222
rect 573 217 589 220
rect 593 223 597 234
rect 601 236 605 241
rect 601 234 602 236
rect 604 234 605 236
rect 601 232 605 234
rect 593 222 616 223
rect 593 220 612 222
rect 614 220 616 222
rect 593 219 616 220
rect 573 215 577 217
rect 572 213 577 215
rect 593 213 597 219
rect 572 211 573 213
rect 575 211 577 213
rect 572 209 577 211
rect 581 212 597 213
rect 581 210 583 212
rect 585 210 597 212
rect 581 209 597 210
rect 500 197 506 198
rect 474 195 489 196
rect 474 193 485 195
rect 487 193 489 195
rect 474 192 489 193
rect 500 195 502 197
rect 504 195 506 197
rect 500 187 506 195
rect 510 197 516 198
rect 510 195 512 197
rect 514 195 516 197
rect 510 194 516 195
rect 573 205 577 209
rect 612 213 616 219
rect 612 209 623 213
rect 573 201 597 205
rect 593 198 597 201
rect 619 203 623 209
rect 619 201 620 203
rect 622 201 623 203
rect 619 199 623 201
rect 593 196 594 198
rect 596 196 597 198
rect 593 194 597 196
rect 604 195 610 196
rect 604 193 606 195
rect 608 193 610 195
rect 533 190 539 191
rect 533 188 535 190
rect 537 188 539 190
rect 533 187 539 188
rect 552 190 558 191
rect 552 188 554 190
rect 556 188 558 190
rect 552 187 558 188
rect 604 187 610 193
rect 17 170 23 171
rect 17 168 19 170
rect 21 168 23 170
rect 17 167 23 168
rect 36 170 42 171
rect 36 168 38 170
rect 40 168 42 170
rect 36 167 42 168
rect 109 165 115 171
rect 71 164 91 165
rect 71 162 87 164
rect 89 162 91 164
rect 109 163 111 165
rect 113 163 115 165
rect 109 162 115 163
rect 122 162 126 164
rect 71 161 91 162
rect 14 157 32 158
rect 14 155 28 157
rect 30 155 32 157
rect 14 154 32 155
rect 14 148 18 154
rect 14 146 15 148
rect 17 146 18 148
rect 10 125 11 136
rect 14 133 18 146
rect 33 141 39 142
rect 59 158 60 160
rect 71 157 75 161
rect 122 160 123 162
rect 125 160 126 162
rect 63 153 75 157
rect 63 148 67 153
rect 63 146 64 148
rect 66 146 67 148
rect 14 129 29 133
rect 25 125 29 129
rect 63 134 67 146
rect 96 157 100 159
rect 96 155 97 157
rect 99 155 100 157
rect 96 149 100 155
rect 122 157 126 160
rect 122 153 146 157
rect 96 145 107 149
rect 63 131 80 134
rect 63 130 77 131
rect 76 129 77 130
rect 79 129 80 131
rect 65 126 71 127
rect 25 124 42 125
rect 25 122 38 124
rect 40 122 42 124
rect 25 121 42 122
rect 65 124 67 126
rect 69 124 71 126
rect 17 117 23 118
rect 17 115 19 117
rect 21 115 23 117
rect 65 115 71 124
rect 76 124 80 129
rect 103 139 107 145
rect 142 149 146 153
rect 122 148 138 149
rect 122 146 134 148
rect 136 146 138 148
rect 122 145 138 146
rect 142 147 147 149
rect 142 145 144 147
rect 146 145 147 147
rect 122 139 126 145
rect 142 143 147 145
rect 142 141 146 143
rect 103 138 126 139
rect 103 136 105 138
rect 107 136 126 138
rect 103 135 126 136
rect 76 122 77 124
rect 79 122 80 124
rect 76 120 80 122
rect 85 124 91 125
rect 85 122 87 124
rect 89 122 91 124
rect 85 115 91 122
rect 114 124 118 126
rect 114 122 115 124
rect 117 122 118 124
rect 114 117 118 122
rect 122 124 126 135
rect 130 138 146 141
rect 130 136 131 138
rect 133 137 146 138
rect 133 136 134 137
rect 130 131 134 136
rect 130 129 131 131
rect 133 129 134 131
rect 130 127 134 129
rect 223 165 229 171
rect 185 164 205 165
rect 185 162 201 164
rect 203 162 205 164
rect 223 163 225 165
rect 227 163 229 165
rect 223 162 229 163
rect 236 162 240 164
rect 185 161 205 162
rect 173 158 174 160
rect 185 157 189 161
rect 236 160 237 162
rect 239 160 240 162
rect 280 164 300 165
rect 280 162 282 164
rect 284 162 300 164
rect 280 161 300 162
rect 177 153 189 157
rect 177 148 181 153
rect 177 146 178 148
rect 180 146 181 148
rect 177 134 181 146
rect 210 157 214 159
rect 210 155 211 157
rect 213 155 214 157
rect 210 149 214 155
rect 236 157 240 160
rect 236 153 260 157
rect 210 145 221 149
rect 177 131 194 134
rect 177 130 191 131
rect 190 129 191 130
rect 193 129 194 131
rect 179 126 185 127
rect 179 124 181 126
rect 183 124 185 126
rect 122 123 155 124
rect 122 121 151 123
rect 153 121 155 123
rect 122 120 155 121
rect 114 115 115 117
rect 117 115 118 117
rect 179 115 185 124
rect 190 124 194 129
rect 217 139 221 145
rect 256 149 260 153
rect 236 148 252 149
rect 236 146 248 148
rect 250 146 252 148
rect 236 145 252 146
rect 256 147 261 149
rect 256 145 258 147
rect 260 145 261 147
rect 236 139 240 145
rect 256 143 261 145
rect 256 141 260 143
rect 217 138 240 139
rect 217 136 219 138
rect 221 136 240 138
rect 217 135 240 136
rect 190 122 191 124
rect 193 122 194 124
rect 190 120 194 122
rect 199 124 205 125
rect 199 122 201 124
rect 203 122 205 124
rect 199 115 205 122
rect 228 124 232 126
rect 228 122 229 124
rect 231 122 232 124
rect 228 117 232 122
rect 236 124 240 135
rect 244 138 260 141
rect 244 136 245 138
rect 247 137 260 138
rect 296 157 300 161
rect 311 158 312 160
rect 296 153 308 157
rect 304 148 308 153
rect 304 146 305 148
rect 307 146 308 148
rect 247 136 248 137
rect 244 131 248 136
rect 244 129 245 131
rect 247 129 248 131
rect 244 127 248 129
rect 304 134 308 146
rect 291 131 308 134
rect 291 129 292 131
rect 294 130 308 131
rect 322 163 328 164
rect 322 161 324 163
rect 326 161 328 163
rect 322 160 328 161
rect 332 163 338 171
rect 332 161 334 163
rect 336 161 338 163
rect 349 165 364 166
rect 349 163 351 165
rect 353 163 364 165
rect 349 162 364 163
rect 332 160 338 161
rect 322 140 326 160
rect 360 157 364 162
rect 367 165 371 171
rect 367 163 368 165
rect 370 163 371 165
rect 367 161 371 163
rect 346 154 357 156
rect 346 152 354 154
rect 356 152 357 154
rect 360 155 374 157
rect 360 153 375 155
rect 346 150 357 152
rect 370 151 372 153
rect 374 151 375 153
rect 346 140 350 150
rect 370 149 375 151
rect 322 139 350 140
rect 322 137 324 139
rect 326 138 350 139
rect 326 137 347 138
rect 322 136 347 137
rect 349 136 350 138
rect 366 139 367 145
rect 346 134 350 136
rect 294 129 295 130
rect 280 124 286 125
rect 236 123 269 124
rect 236 121 265 123
rect 267 121 269 123
rect 236 120 269 121
rect 280 122 282 124
rect 284 122 286 124
rect 228 115 229 117
rect 231 115 232 117
rect 280 115 286 122
rect 291 124 295 129
rect 370 132 374 149
rect 358 128 374 132
rect 291 122 292 124
rect 294 122 295 124
rect 291 120 295 122
rect 300 126 306 127
rect 300 124 302 126
rect 304 124 306 126
rect 300 115 306 124
rect 349 127 362 128
rect 349 125 351 127
rect 353 125 362 127
rect 349 124 362 125
rect 400 165 404 171
rect 400 163 401 165
rect 403 163 404 165
rect 400 161 404 163
rect 407 165 422 166
rect 407 163 418 165
rect 420 163 422 165
rect 407 162 422 163
rect 433 163 439 171
rect 467 165 471 171
rect 407 157 411 162
rect 433 161 435 163
rect 437 161 439 163
rect 433 160 439 161
rect 443 163 449 164
rect 443 161 445 163
rect 447 161 449 163
rect 443 160 449 161
rect 397 155 411 157
rect 396 153 411 155
rect 414 154 425 156
rect 396 151 397 153
rect 399 151 401 153
rect 396 149 401 151
rect 414 152 415 154
rect 417 152 425 154
rect 414 150 425 152
rect 397 132 401 149
rect 404 139 405 145
rect 421 140 425 150
rect 445 140 449 160
rect 421 139 449 140
rect 421 138 445 139
rect 421 136 422 138
rect 424 137 445 138
rect 447 137 449 139
rect 424 136 449 137
rect 467 163 468 165
rect 470 163 471 165
rect 467 161 471 163
rect 474 165 489 166
rect 474 163 485 165
rect 487 163 489 165
rect 474 162 489 163
rect 500 163 506 171
rect 533 170 539 171
rect 533 168 535 170
rect 537 168 539 170
rect 533 167 539 168
rect 552 170 558 171
rect 552 168 554 170
rect 556 168 558 170
rect 552 167 558 168
rect 604 165 610 171
rect 474 157 478 162
rect 500 161 502 163
rect 504 161 506 163
rect 500 160 506 161
rect 510 163 516 164
rect 510 161 512 163
rect 514 161 516 163
rect 510 160 516 161
rect 464 155 478 157
rect 421 134 425 136
rect 397 128 413 132
rect 409 127 422 128
rect 409 125 418 127
rect 420 125 422 127
rect 409 124 422 125
rect 463 153 478 155
rect 481 154 492 156
rect 463 151 464 153
rect 466 151 468 153
rect 463 149 468 151
rect 481 152 482 154
rect 484 152 492 154
rect 481 150 492 152
rect 464 132 468 149
rect 471 139 472 145
rect 488 140 492 150
rect 512 140 516 160
rect 593 162 597 164
rect 604 163 606 165
rect 608 163 610 165
rect 604 162 610 163
rect 488 139 516 140
rect 488 138 512 139
rect 488 136 489 138
rect 491 137 512 138
rect 514 137 516 139
rect 491 136 516 137
rect 530 157 548 158
rect 530 155 544 157
rect 546 155 548 157
rect 530 154 548 155
rect 488 134 492 136
rect 530 148 534 154
rect 530 146 531 148
rect 533 146 534 148
rect 464 128 480 132
rect 476 127 489 128
rect 476 125 485 127
rect 487 125 489 127
rect 476 124 489 125
rect 526 125 527 136
rect 530 133 534 146
rect 593 160 594 162
rect 596 160 597 162
rect 593 157 597 160
rect 549 141 555 142
rect 530 129 545 133
rect 541 125 545 129
rect 573 153 597 157
rect 573 149 577 153
rect 619 157 623 159
rect 619 155 620 157
rect 622 155 623 157
rect 572 147 577 149
rect 572 145 573 147
rect 575 145 577 147
rect 581 148 597 149
rect 581 146 583 148
rect 585 146 597 148
rect 581 145 597 146
rect 572 143 577 145
rect 573 141 577 143
rect 573 138 589 141
rect 573 137 586 138
rect 585 136 586 137
rect 588 136 589 138
rect 585 131 589 136
rect 585 129 586 131
rect 588 129 589 131
rect 585 127 589 129
rect 593 139 597 145
rect 619 149 623 155
rect 612 145 623 149
rect 612 139 616 145
rect 593 138 616 139
rect 593 136 612 138
rect 614 136 616 138
rect 593 135 616 136
rect 541 124 558 125
rect 593 124 597 135
rect 541 122 554 124
rect 556 122 558 124
rect 541 121 558 122
rect 564 123 597 124
rect 564 121 566 123
rect 568 121 597 123
rect 564 120 597 121
rect 601 124 605 126
rect 601 122 602 124
rect 604 122 605 124
rect 333 117 337 119
rect 333 115 334 117
rect 336 115 337 117
rect 366 117 372 118
rect 366 115 368 117
rect 370 115 372 117
rect 399 117 405 118
rect 399 115 401 117
rect 403 115 405 117
rect 434 117 438 119
rect 434 115 435 117
rect 437 115 438 117
rect 466 117 472 118
rect 466 115 468 117
rect 470 115 472 117
rect 501 117 505 119
rect 501 115 502 117
rect 504 115 505 117
rect 533 117 539 118
rect 533 115 535 117
rect 537 115 539 117
rect 601 117 605 122
rect 601 115 602 117
rect 604 115 605 117
rect 17 97 19 99
rect 21 97 23 99
rect 17 96 23 97
rect 25 92 42 93
rect 25 90 38 92
rect 40 90 42 92
rect 25 89 42 90
rect 65 90 71 99
rect 10 78 11 89
rect 25 85 29 89
rect 65 88 67 90
rect 69 88 71 90
rect 65 87 71 88
rect 76 92 80 94
rect 76 90 77 92
rect 79 90 80 92
rect 14 81 29 85
rect 76 85 80 90
rect 85 92 91 99
rect 114 97 115 99
rect 117 97 118 99
rect 85 90 87 92
rect 89 90 91 92
rect 85 89 91 90
rect 114 92 118 97
rect 114 90 115 92
rect 117 90 118 92
rect 114 88 118 90
rect 122 93 155 94
rect 122 91 151 93
rect 153 91 155 93
rect 122 90 155 91
rect 179 90 185 99
rect 76 84 77 85
rect 14 68 18 81
rect 63 83 77 84
rect 79 83 80 85
rect 63 80 80 83
rect 33 72 39 73
rect 14 66 15 68
rect 17 66 18 68
rect 14 60 18 66
rect 14 59 32 60
rect 14 57 28 59
rect 30 57 32 59
rect 14 56 32 57
rect 63 68 67 80
rect 122 79 126 90
rect 179 88 181 90
rect 183 88 185 90
rect 179 87 185 88
rect 190 92 194 94
rect 190 90 191 92
rect 193 90 194 92
rect 103 78 126 79
rect 103 76 105 78
rect 107 76 126 78
rect 103 75 126 76
rect 103 69 107 75
rect 63 66 64 68
rect 66 66 67 68
rect 63 61 67 66
rect 63 57 75 61
rect 59 54 60 56
rect 71 53 75 57
rect 96 65 107 69
rect 96 59 100 65
rect 122 69 126 75
rect 130 85 134 87
rect 130 83 131 85
rect 133 83 134 85
rect 130 78 134 83
rect 130 76 131 78
rect 133 77 134 78
rect 133 76 146 77
rect 130 73 146 76
rect 142 71 146 73
rect 142 69 147 71
rect 122 68 138 69
rect 122 66 134 68
rect 136 66 138 68
rect 122 65 138 66
rect 142 67 144 69
rect 146 67 147 69
rect 142 65 147 67
rect 96 57 97 59
rect 99 57 100 59
rect 96 55 100 57
rect 142 61 146 65
rect 122 57 146 61
rect 122 54 126 57
rect 71 52 91 53
rect 122 52 123 54
rect 125 52 126 54
rect 71 50 87 52
rect 89 50 91 52
rect 71 49 91 50
rect 109 51 115 52
rect 109 49 111 51
rect 113 49 115 51
rect 122 50 126 52
rect 190 85 194 90
rect 199 92 205 99
rect 228 97 229 99
rect 231 97 232 99
rect 199 90 201 92
rect 203 90 205 92
rect 199 89 205 90
rect 228 92 232 97
rect 228 90 229 92
rect 231 90 232 92
rect 228 88 232 90
rect 236 93 269 94
rect 236 91 265 93
rect 267 91 269 93
rect 236 90 269 91
rect 280 92 286 99
rect 280 90 282 92
rect 284 90 286 92
rect 190 84 191 85
rect 177 83 191 84
rect 193 83 194 85
rect 177 80 194 83
rect 177 68 181 80
rect 236 79 240 90
rect 280 89 286 90
rect 291 92 295 94
rect 291 90 292 92
rect 294 90 295 92
rect 217 78 240 79
rect 217 76 219 78
rect 221 76 240 78
rect 217 75 240 76
rect 217 69 221 75
rect 177 66 178 68
rect 180 66 181 68
rect 177 61 181 66
rect 177 57 189 61
rect 173 54 174 56
rect 17 46 23 47
rect 17 44 19 46
rect 21 44 23 46
rect 17 43 23 44
rect 36 46 42 47
rect 36 44 38 46
rect 40 44 42 46
rect 36 43 42 44
rect 109 43 115 49
rect 185 53 189 57
rect 210 65 221 69
rect 210 59 214 65
rect 236 69 240 75
rect 244 85 248 87
rect 244 83 245 85
rect 247 83 248 85
rect 244 78 248 83
rect 244 76 245 78
rect 247 77 248 78
rect 247 76 260 77
rect 244 73 260 76
rect 256 71 260 73
rect 291 85 295 90
rect 300 90 306 99
rect 333 97 334 99
rect 336 97 337 99
rect 333 95 337 97
rect 366 97 368 99
rect 370 97 372 99
rect 366 96 372 97
rect 399 97 401 99
rect 403 97 405 99
rect 399 96 405 97
rect 434 97 435 99
rect 437 97 438 99
rect 434 95 438 97
rect 466 97 468 99
rect 470 97 472 99
rect 466 96 472 97
rect 501 97 502 99
rect 504 97 505 99
rect 501 95 505 97
rect 533 97 535 99
rect 537 97 539 99
rect 533 96 539 97
rect 601 97 602 99
rect 604 97 605 99
rect 300 88 302 90
rect 304 88 306 90
rect 300 87 306 88
rect 291 83 292 85
rect 294 84 295 85
rect 294 83 308 84
rect 291 80 308 83
rect 256 69 261 71
rect 236 68 252 69
rect 236 66 248 68
rect 250 66 252 68
rect 236 65 252 66
rect 256 67 258 69
rect 260 67 261 69
rect 256 65 261 67
rect 210 57 211 59
rect 213 57 214 59
rect 210 55 214 57
rect 256 61 260 65
rect 236 57 260 61
rect 236 54 240 57
rect 185 52 205 53
rect 236 52 237 54
rect 239 52 240 54
rect 304 68 308 80
rect 349 89 362 90
rect 349 87 351 89
rect 353 87 362 89
rect 349 86 362 87
rect 358 82 374 86
rect 346 78 350 80
rect 304 66 305 68
rect 307 66 308 68
rect 304 61 308 66
rect 296 57 308 61
rect 296 53 300 57
rect 311 54 312 56
rect 185 50 201 52
rect 203 50 205 52
rect 185 49 205 50
rect 223 51 229 52
rect 223 49 225 51
rect 227 49 229 51
rect 236 50 240 52
rect 280 52 300 53
rect 280 50 282 52
rect 284 50 300 52
rect 280 49 300 50
rect 223 43 229 49
rect 322 77 347 78
rect 322 75 324 77
rect 326 76 347 77
rect 349 76 350 78
rect 326 75 350 76
rect 322 74 350 75
rect 322 54 326 74
rect 346 64 350 74
rect 366 69 367 75
rect 370 65 374 82
rect 346 62 357 64
rect 346 60 354 62
rect 356 60 357 62
rect 370 63 375 65
rect 370 61 372 63
rect 374 61 375 63
rect 346 58 357 60
rect 360 59 375 61
rect 360 57 374 59
rect 322 53 328 54
rect 322 51 324 53
rect 326 51 328 53
rect 322 50 328 51
rect 332 53 338 54
rect 332 51 334 53
rect 336 51 338 53
rect 360 52 364 57
rect 332 43 338 51
rect 349 51 364 52
rect 349 49 351 51
rect 353 49 364 51
rect 349 48 364 49
rect 367 51 371 53
rect 367 49 368 51
rect 370 49 371 51
rect 367 43 371 49
rect 409 89 422 90
rect 409 87 418 89
rect 420 87 422 89
rect 409 86 422 87
rect 397 82 413 86
rect 397 65 401 82
rect 476 89 489 90
rect 421 78 425 80
rect 404 69 405 75
rect 421 76 422 78
rect 424 77 449 78
rect 424 76 445 77
rect 421 75 445 76
rect 447 75 449 77
rect 421 74 449 75
rect 396 63 401 65
rect 421 64 425 74
rect 396 61 397 63
rect 399 61 401 63
rect 414 62 425 64
rect 396 59 411 61
rect 397 57 411 59
rect 414 60 415 62
rect 417 60 425 62
rect 414 58 425 60
rect 400 51 404 53
rect 400 49 401 51
rect 403 49 404 51
rect 400 43 404 49
rect 407 52 411 57
rect 445 54 449 74
rect 433 53 439 54
rect 407 51 422 52
rect 407 49 418 51
rect 420 49 422 51
rect 407 48 422 49
rect 433 51 435 53
rect 437 51 439 53
rect 433 43 439 51
rect 443 53 449 54
rect 443 51 445 53
rect 447 51 449 53
rect 443 50 449 51
rect 476 87 485 89
rect 487 87 489 89
rect 476 86 489 87
rect 464 82 480 86
rect 464 65 468 82
rect 564 93 597 94
rect 541 92 558 93
rect 541 90 554 92
rect 556 90 558 92
rect 564 91 566 93
rect 568 91 597 93
rect 564 90 597 91
rect 541 89 558 90
rect 488 78 492 80
rect 471 69 472 75
rect 488 76 489 78
rect 491 77 516 78
rect 491 76 512 77
rect 488 75 512 76
rect 514 75 516 77
rect 488 74 516 75
rect 463 63 468 65
rect 488 64 492 74
rect 463 61 464 63
rect 466 61 468 63
rect 481 62 492 64
rect 463 59 478 61
rect 464 57 478 59
rect 481 60 482 62
rect 484 60 492 62
rect 481 58 492 60
rect 467 51 471 53
rect 467 49 468 51
rect 470 49 471 51
rect 467 43 471 49
rect 474 52 478 57
rect 512 54 516 74
rect 526 78 527 89
rect 541 85 545 89
rect 530 81 545 85
rect 530 68 534 81
rect 585 85 589 87
rect 585 83 586 85
rect 588 83 589 85
rect 549 72 555 73
rect 530 66 531 68
rect 533 66 534 68
rect 530 60 534 66
rect 530 59 548 60
rect 530 57 544 59
rect 546 57 548 59
rect 530 56 548 57
rect 585 78 589 83
rect 585 77 586 78
rect 573 76 586 77
rect 588 76 589 78
rect 573 73 589 76
rect 593 79 597 90
rect 601 92 605 97
rect 601 90 602 92
rect 604 90 605 92
rect 601 88 605 90
rect 593 78 616 79
rect 593 76 612 78
rect 614 76 616 78
rect 593 75 616 76
rect 573 71 577 73
rect 572 69 577 71
rect 593 69 597 75
rect 572 67 573 69
rect 575 67 577 69
rect 572 65 577 67
rect 581 68 597 69
rect 581 66 583 68
rect 585 66 597 68
rect 581 65 597 66
rect 500 53 506 54
rect 474 51 489 52
rect 474 49 485 51
rect 487 49 489 51
rect 474 48 489 49
rect 500 51 502 53
rect 504 51 506 53
rect 500 43 506 51
rect 510 53 516 54
rect 510 51 512 53
rect 514 51 516 53
rect 510 50 516 51
rect 573 61 577 65
rect 612 69 616 75
rect 612 65 623 69
rect 573 57 597 61
rect 593 54 597 57
rect 619 59 623 65
rect 619 57 620 59
rect 622 57 623 59
rect 619 55 623 57
rect 593 52 594 54
rect 596 52 597 54
rect 593 50 597 52
rect 604 51 610 52
rect 604 49 606 51
rect 608 49 610 51
rect 533 46 539 47
rect 533 44 535 46
rect 537 44 539 46
rect 533 43 539 44
rect 552 46 558 47
rect 552 44 554 46
rect 556 44 558 46
rect 552 43 558 44
rect 604 43 610 49
<< via1 >>
rect 39 290 41 292
rect 80 299 82 301
rect 105 299 107 301
rect 88 275 90 277
rect 152 298 154 300
rect 97 275 99 277
rect 170 290 172 292
rect 194 299 196 301
rect 219 299 221 301
rect 202 275 204 277
rect 211 275 213 277
rect 266 283 268 285
rect 313 298 315 300
rect 330 298 332 300
rect 355 282 357 284
rect 332 274 334 276
rect 379 290 381 292
rect 406 290 408 292
rect 437 298 439 300
rect 457 298 459 300
rect 480 283 482 285
rect 505 298 507 300
rect 523 282 525 284
rect 504 274 506 276
rect 565 298 567 300
rect 7 219 9 221
rect 88 225 90 227
rect 39 210 41 212
rect 97 225 99 227
rect 80 201 82 203
rect 105 201 107 203
rect 152 202 154 204
rect 202 225 204 227
rect 170 210 172 212
rect 211 225 213 227
rect 194 201 196 203
rect 266 217 268 219
rect 219 201 221 203
rect 332 226 334 228
rect 313 202 315 204
rect 330 202 332 204
rect 355 218 357 220
rect 379 210 381 212
rect 406 210 408 212
rect 437 202 439 204
rect 504 226 506 228
rect 480 217 482 219
rect 457 202 459 204
rect 505 202 507 204
rect 523 218 525 220
rect 565 202 567 204
rect 7 147 9 149
rect 39 146 41 148
rect 80 155 82 157
rect 105 155 107 157
rect 88 131 90 133
rect 152 154 154 156
rect 97 131 99 133
rect 170 146 172 148
rect 194 155 196 157
rect 219 155 221 157
rect 202 131 204 133
rect 211 131 213 133
rect 266 139 268 141
rect 313 154 315 156
rect 330 154 332 156
rect 355 138 357 140
rect 332 130 334 132
rect 379 146 381 148
rect 406 146 408 148
rect 437 154 439 156
rect 457 154 459 156
rect 480 139 482 141
rect 505 154 507 156
rect 523 138 525 140
rect 504 130 506 132
rect 565 154 567 156
rect 7 75 9 77
rect 88 81 90 83
rect 39 66 41 68
rect 97 81 99 83
rect 80 57 82 59
rect 105 57 107 59
rect 152 58 154 60
rect 202 81 204 83
rect 170 66 172 68
rect 211 81 213 83
rect 194 57 196 59
rect 266 73 268 75
rect 219 57 221 59
rect 332 82 334 84
rect 313 58 315 60
rect 330 58 332 60
rect 355 74 357 76
rect 379 66 381 68
rect 406 66 408 68
rect 437 58 439 60
rect 504 82 506 84
rect 480 73 482 75
rect 457 58 459 60
rect 505 58 507 60
rect 523 74 525 76
rect 565 58 567 60
<< labels >>
rlabel alu1 125 319 125 319 8 vss
rlabel alu1 125 255 125 255 8 vdd
rlabel alu1 73 255 73 255 8 vdd
rlabel alu1 73 319 73 319 8 vss
rlabel alu1 239 319 239 319 8 vss
rlabel alu1 239 255 239 255 8 vdd
rlabel alu1 267 295 267 295 5 sum
rlabel alu1 187 255 187 255 8 vdd
rlabel alu1 187 319 187 319 8 vss
rlabel alu1 24 319 24 319 8 vss
rlabel alu1 24 255 24 255 8 vdd
rlabel alu1 298 319 298 319 2 vss
rlabel alu1 298 255 298 255 2 vdd
rlabel alu1 419 319 419 319 8 vss
rlabel alu1 419 255 419 255 8 vdd
rlabel alu1 352 319 352 319 2 vss
rlabel alu1 352 255 352 255 2 vdd
rlabel alu1 486 319 486 319 8 vss
rlabel alu1 486 255 486 255 8 vdd
rlabel via1 506 275 506 275 5 s1
rlabel alu1 514 267 514 267 5 s1
rlabel via1 332 275 332 275 5 s1
rlabel alu1 324 267 324 267 5 s1
rlabel alu1 447 267 447 267 5 s0
rlabel alu1 540 319 540 319 8 vss
rlabel alu1 540 255 540 255 8 vdd
rlabel alu1 594 319 594 319 2 vss
rlabel alu1 594 255 594 255 2 vdd
rlabel via1 332 299 332 299 1 i1
rlabel via1 356 283 356 283 1 i0
rlabel alu1 340 291 340 291 1 i1
rlabel polyct1 364 287 364 287 1 i0
rlabel alu1 474 289 474 289 1 i2
rlabel alu1 478 284 478 284 1 i2
rlabel alu1 497 291 497 291 1 i3
rlabel alu1 502 300 502 300 1 i3
rlabel alu1 8 289 8 289 1 cout3
rlabel alu2 73 292 73 292 1 a3
rlabel via1 88 277 88 277 1 b3
rlabel alu1 290 295 290 295 1 a3
rlabel alu1 298 291 298 291 1 a3
rlabel alu2 290 283 290 283 1 b3
rlabel alu1 282 275 282 275 1 b3
rlabel alu1 391 286 391 286 1 z3
rlabel alu1 399 267 399 267 1 z3
rlabel alu1 540 291 540 291 1 a3
rlabel alu1 548 291 548 291 1 a3
rlabel alu2 556 299 556 299 1 a3
rlabel alu1 540 283 540 283 1 b3
rlabel alu1 548 283 548 283 1 b3
rlabel alu1 556 275 556 275 1 b3
rlabel polyct1 606 295 606 295 1 a3
rlabel alu1 614 299 614 299 1 a3
rlabel alu1 622 275 622 275 1 b3
rlabel alu1 614 267 614 267 1 b3
rlabel alu1 125 183 125 183 6 vss
rlabel alu1 125 247 125 247 6 vdd
rlabel alu1 73 247 73 247 6 vdd
rlabel alu1 73 183 73 183 6 vss
rlabel alu1 239 183 239 183 6 vss
rlabel alu1 239 247 239 247 6 vdd
rlabel alu1 267 207 267 207 1 sum
rlabel alu1 187 247 187 247 6 vdd
rlabel alu1 187 183 187 183 6 vss
rlabel alu1 24 183 24 183 6 vss
rlabel alu1 24 247 24 247 6 vdd
rlabel alu1 298 183 298 183 4 vss
rlabel alu1 298 247 298 247 4 vdd
rlabel alu1 419 183 419 183 6 vss
rlabel alu1 419 247 419 247 6 vdd
rlabel alu1 352 183 352 183 4 vss
rlabel alu1 352 247 352 247 4 vdd
rlabel alu1 486 183 486 183 6 vss
rlabel alu1 486 247 486 247 6 vdd
rlabel via1 506 227 506 227 1 s1
rlabel alu1 514 235 514 235 1 s1
rlabel via1 332 227 332 227 1 s1
rlabel alu1 324 235 324 235 1 s1
rlabel alu1 447 235 447 235 1 s0
rlabel alu1 540 183 540 183 6 vss
rlabel alu1 540 247 540 247 6 vdd
rlabel alu1 594 183 594 183 4 vss
rlabel alu1 594 247 594 247 4 vdd
rlabel via1 332 203 332 203 1 i1
rlabel alu1 340 211 340 211 1 i1
rlabel via1 356 219 356 219 1 i0
rlabel polyct1 364 215 364 215 1 i1
rlabel alu1 474 213 474 213 1 i2
rlabel alu1 478 218 478 218 1 i2
rlabel alu1 497 211 497 211 1 i3
rlabel alu1 502 202 502 202 1 i3
rlabel alu1 8 213 8 213 1 cout2
rlabel alu2 73 210 73 210 1 a2
rlabel via1 88 225 88 225 1 a2
rlabel alu1 282 227 282 227 1 b2
rlabel alu2 290 219 290 219 1 b2
rlabel alu1 290 207 290 207 1 a2
rlabel alu1 298 211 298 211 1 a2
rlabel alu1 540 219 540 219 1 b2
rlabel alu1 548 219 548 219 1 b2
rlabel alu1 556 227 556 227 1 b2
rlabel alu1 540 211 540 211 1 a2
rlabel alu1 548 211 548 211 1 a2
rlabel alu1 614 235 614 235 1 b2
rlabel alu1 622 227 622 227 1 b2
rlabel polyct1 606 207 606 207 1 a2
rlabel alu1 614 203 614 203 1 a2
rlabel alu1 391 216 391 216 1 z2
rlabel alu1 399 235 399 235 1 z2
rlabel alu2 8 145 8 145 1 cout1
rlabel alu1 391 142 391 142 1 z1
rlabel alu1 614 155 614 155 1 a1
rlabel polyct1 606 151 606 151 1 a1
rlabel alu1 622 131 622 131 1 b1
rlabel alu1 614 123 614 123 1 b1
rlabel alu1 556 131 556 131 1 b1
rlabel alu1 548 139 548 139 1 b1
rlabel alu1 540 139 540 139 1 b1
rlabel alu2 556 155 556 155 1 a1
rlabel alu1 548 147 548 147 1 a1
rlabel alu1 540 147 540 147 1 a1
rlabel alu1 502 156 502 156 1 i3
rlabel alu1 497 147 497 147 1 i3
rlabel alu1 478 140 478 140 1 i2
rlabel alu1 474 145 474 145 1 i2
rlabel alu1 399 123 399 123 1 z1
rlabel polyct1 364 143 364 143 1 i0
rlabel alu1 340 147 340 147 1 i1
rlabel via1 356 139 356 139 1 i0
rlabel via1 332 155 332 155 1 i1
rlabel alu1 282 131 282 131 1 b1
rlabel alu2 290 139 290 139 1 b1
rlabel alu1 298 147 298 147 1 a1
rlabel alu1 290 151 290 151 1 a1
rlabel via1 88 133 88 133 1 b1
rlabel alu2 73 148 73 148 1 a1
rlabel alu1 594 111 594 111 2 vdd
rlabel alu1 594 175 594 175 2 vss
rlabel alu1 540 111 540 111 8 vdd
rlabel alu1 540 175 540 175 8 vss
rlabel alu1 447 123 447 123 5 s0
rlabel alu1 324 123 324 123 5 s1
rlabel via1 332 131 332 131 5 s1
rlabel alu1 514 123 514 123 5 s1
rlabel via1 506 131 506 131 5 s1
rlabel alu1 486 111 486 111 8 vdd
rlabel alu1 486 175 486 175 8 vss
rlabel alu1 352 111 352 111 2 vdd
rlabel alu1 352 175 352 175 2 vss
rlabel alu1 419 111 419 111 8 vdd
rlabel alu1 419 175 419 175 8 vss
rlabel alu1 298 111 298 111 2 vdd
rlabel alu1 298 175 298 175 2 vss
rlabel alu1 24 111 24 111 8 vdd
rlabel alu1 24 175 24 175 8 vss
rlabel alu1 187 175 187 175 8 vss
rlabel alu1 187 111 187 111 8 vdd
rlabel alu1 267 151 267 151 5 sum
rlabel alu1 239 111 239 111 8 vdd
rlabel alu1 239 175 239 175 8 vss
rlabel alu1 73 175 73 175 8 vss
rlabel alu1 73 111 73 111 8 vdd
rlabel alu1 125 111 125 111 8 vdd
rlabel alu1 125 175 125 175 8 vss
rlabel alu1 8 69 8 69 1 cout0
rlabel alu1 399 91 399 91 1 z0
rlabel alu1 622 83 622 83 1 b0
rlabel alu1 614 91 614 91 1 b0
rlabel alu1 614 59 614 59 1 a0
rlabel polyct1 606 63 606 63 1 a0
rlabel alu1 556 83 556 83 1 b0
rlabel alu1 548 75 548 75 1 b0
rlabel alu1 540 75 540 75 1 b0
rlabel alu1 540 67 540 67 1 a0
rlabel alu1 548 67 548 67 1 a0
rlabel alu1 502 58 502 58 1 i3
rlabel alu1 497 67 497 67 1 i3
rlabel alu1 478 74 478 74 1 i2
rlabel alu1 474 69 474 69 1 i2
rlabel alu1 391 72 391 72 1 z0
rlabel polyct1 364 71 364 71 1 i1
rlabel via1 356 75 356 75 1 i0
rlabel alu1 340 67 340 67 1 i1
rlabel via1 332 59 332 59 1 i1
rlabel alu2 290 75 290 75 1 b0
rlabel alu1 282 83 282 83 1 b0
rlabel alu1 298 67 298 67 1 a0
rlabel alu1 290 63 290 63 1 a0
rlabel via1 88 81 88 81 1 b0
rlabel alu2 73 66 73 66 1 a0
rlabel alu1 594 103 594 103 4 vdd
rlabel alu1 594 39 594 39 4 vss
rlabel alu1 540 103 540 103 6 vdd
rlabel alu1 540 39 540 39 6 vss
rlabel alu1 447 91 447 91 1 s0
rlabel alu1 324 91 324 91 1 s1
rlabel via1 332 83 332 83 1 s1
rlabel alu1 514 91 514 91 1 s1
rlabel via1 506 83 506 83 1 s1
rlabel alu1 486 103 486 103 6 vdd
rlabel alu1 486 39 486 39 6 vss
rlabel alu1 352 103 352 103 4 vdd
rlabel alu1 352 39 352 39 4 vss
rlabel alu1 419 103 419 103 6 vdd
rlabel alu1 419 39 419 39 6 vss
rlabel alu1 298 103 298 103 4 vdd
rlabel alu1 298 39 298 39 4 vss
rlabel via1 204 82 204 82 1 cin
rlabel alu1 24 103 24 103 6 vdd
rlabel alu1 24 39 24 39 6 vss
rlabel alu1 187 39 187 39 6 vss
rlabel alu1 187 103 187 103 6 vdd
rlabel alu1 267 63 267 63 1 sum
rlabel alu1 239 103 239 103 6 vdd
rlabel alu1 239 39 239 39 6 vss
rlabel alu1 73 39 73 39 6 vss
rlabel alu1 73 103 73 103 6 vdd
rlabel alu1 125 103 125 103 6 vdd
rlabel alu1 125 39 125 39 6 vss
<< end >>
