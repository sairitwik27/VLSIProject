magic
tech scmos
timestamp 1607760857
<< ab >>
rect 84 148 90 153
rect 198 148 204 153
rect 0 76 40 148
rect 49 116 153 148
rect 49 84 89 116
rect 90 84 153 116
rect 42 76 47 84
rect 49 76 153 84
rect 163 116 267 148
rect 268 140 272 148
rect 163 84 203 116
rect 204 84 267 116
rect 163 76 267 84
rect 268 76 270 84
rect 274 76 314 148
rect 315 140 379 148
rect 318 84 379 140
rect 315 76 379 84
rect 383 76 447 148
rect 451 76 514 148
rect 516 140 556 148
rect 558 140 628 148
rect 517 84 556 140
rect 559 84 622 140
rect 516 76 556 84
rect 557 76 622 84
rect 623 76 628 84
rect 1 4 41 76
rect 43 68 48 76
rect 50 68 154 76
rect 50 36 90 68
rect 91 36 154 68
rect 50 4 154 36
rect 164 68 268 76
rect 269 68 271 76
rect 164 36 204 68
rect 205 36 268 68
rect 164 4 268 36
rect 269 4 273 12
rect 275 4 315 76
rect 316 68 380 76
rect 319 12 380 68
rect 316 4 380 12
rect 384 4 448 76
rect 452 4 515 76
rect 517 68 557 76
rect 558 68 623 76
rect 624 68 629 76
rect 518 12 557 68
rect 560 12 623 68
rect 517 4 557 12
rect 559 4 629 12
rect 85 -1 91 4
rect 199 -1 205 4
<< nwell >>
rect -5 81 628 116
rect -5 71 629 81
rect -4 36 629 71
<< pwell >>
rect -5 116 628 153
rect -4 -1 629 36
<< poly >>
rect 9 131 11 136
rect 19 128 21 133
rect 29 128 31 133
rect 58 133 60 137
rect 71 135 73 140
rect 78 135 80 140
rect 101 144 126 146
rect 101 136 103 144
rect 114 136 116 140
rect 124 136 126 144
rect 134 139 136 144
rect 141 139 143 144
rect 98 134 103 136
rect 98 131 100 134
rect 9 119 11 122
rect 19 119 21 122
rect 9 117 15 119
rect 9 115 11 117
rect 13 115 15 117
rect 9 113 15 115
rect 19 117 25 119
rect 19 115 21 117
rect 23 115 25 117
rect 19 113 25 115
rect 9 110 11 113
rect 22 103 24 113
rect 29 112 31 122
rect 58 119 60 124
rect 71 119 73 124
rect 58 117 64 119
rect 58 115 60 117
rect 62 115 64 117
rect 58 113 64 115
rect 68 117 74 119
rect 68 115 70 117
rect 72 115 74 117
rect 68 113 74 115
rect 29 110 35 112
rect 29 108 31 110
rect 33 108 35 110
rect 58 109 60 113
rect 29 106 35 108
rect 29 103 31 106
rect 9 87 11 92
rect 68 102 70 113
rect 78 111 80 124
rect 172 133 174 137
rect 185 135 187 140
rect 192 135 194 140
rect 215 144 240 146
rect 215 136 217 144
rect 228 136 230 140
rect 238 136 240 144
rect 248 139 250 144
rect 255 139 257 144
rect 114 124 116 127
rect 107 122 116 124
rect 124 123 126 127
rect 134 124 136 127
rect 98 114 100 122
rect 107 120 109 122
rect 111 120 116 122
rect 107 118 116 120
rect 132 122 136 124
rect 132 119 134 122
rect 114 114 116 118
rect 128 117 134 119
rect 141 118 143 127
rect 212 134 217 136
rect 212 131 214 134
rect 172 119 174 124
rect 185 119 187 124
rect 128 115 130 117
rect 132 115 134 117
rect 95 112 108 114
rect 114 112 124 114
rect 128 113 134 115
rect 95 111 97 112
rect 78 109 84 111
rect 78 107 80 109
rect 82 107 84 109
rect 78 105 84 107
rect 91 109 97 111
rect 106 109 108 112
rect 122 109 124 112
rect 132 109 134 113
rect 138 116 144 118
rect 138 114 140 116
rect 142 114 144 116
rect 138 112 144 114
rect 142 109 144 112
rect 172 117 178 119
rect 172 115 174 117
rect 176 115 178 117
rect 172 113 178 115
rect 182 117 188 119
rect 182 115 184 117
rect 186 115 188 117
rect 182 113 188 115
rect 172 109 174 113
rect 91 107 93 109
rect 95 107 97 109
rect 91 105 97 107
rect 78 102 80 105
rect 58 87 60 91
rect 68 84 70 89
rect 78 84 80 89
rect 22 78 24 82
rect 29 78 31 82
rect 122 87 124 91
rect 132 87 134 91
rect 106 78 108 82
rect 182 102 184 113
rect 192 111 194 124
rect 283 135 285 140
rect 290 135 292 140
rect 325 144 344 146
rect 228 124 230 127
rect 221 122 230 124
rect 238 123 240 127
rect 248 124 250 127
rect 212 114 214 122
rect 221 120 223 122
rect 225 120 230 122
rect 221 118 230 120
rect 246 122 250 124
rect 246 119 248 122
rect 228 114 230 118
rect 242 117 248 119
rect 255 118 257 127
rect 303 133 305 137
rect 325 134 327 144
rect 335 136 337 140
rect 342 136 344 144
rect 419 144 438 146
rect 352 136 354 141
rect 359 136 361 141
rect 369 136 371 141
rect 392 136 394 141
rect 402 136 404 141
rect 409 136 411 141
rect 419 136 421 144
rect 426 136 428 140
rect 242 115 244 117
rect 246 115 248 117
rect 209 112 222 114
rect 228 112 238 114
rect 242 113 248 115
rect 209 111 211 112
rect 192 109 198 111
rect 192 107 194 109
rect 196 107 198 109
rect 192 105 198 107
rect 205 109 211 111
rect 220 109 222 112
rect 236 109 238 112
rect 246 109 248 113
rect 252 116 258 118
rect 252 114 254 116
rect 256 114 258 116
rect 252 112 258 114
rect 256 109 258 112
rect 283 111 285 124
rect 290 119 292 124
rect 303 119 305 124
rect 289 117 295 119
rect 289 115 291 117
rect 293 115 295 117
rect 289 113 295 115
rect 299 117 305 119
rect 299 115 301 117
rect 303 115 305 117
rect 299 113 305 115
rect 279 109 285 111
rect 205 107 207 109
rect 209 107 211 109
rect 205 105 211 107
rect 192 102 194 105
rect 172 87 174 91
rect 182 84 184 89
rect 192 84 194 89
rect 142 78 144 82
rect 236 87 238 91
rect 246 87 248 91
rect 220 78 222 82
rect 279 107 281 109
rect 283 107 285 109
rect 279 105 285 107
rect 283 102 285 105
rect 293 102 295 113
rect 303 109 305 113
rect 325 110 327 128
rect 335 119 337 128
rect 331 117 337 119
rect 331 115 333 117
rect 335 115 337 117
rect 331 113 337 115
rect 342 115 344 128
rect 352 125 354 128
rect 348 123 354 125
rect 348 121 350 123
rect 352 121 354 123
rect 348 119 354 121
rect 342 113 354 115
rect 359 114 361 128
rect 436 134 438 144
rect 486 144 505 146
rect 459 136 461 141
rect 469 136 471 141
rect 476 136 478 141
rect 486 136 488 144
rect 493 136 495 140
rect 369 124 371 127
rect 392 124 394 127
rect 366 122 372 124
rect 366 120 368 122
rect 370 120 372 122
rect 366 118 372 120
rect 391 122 397 124
rect 391 120 393 122
rect 395 120 397 122
rect 391 118 397 120
rect 325 99 327 102
rect 318 97 327 99
rect 335 98 337 113
rect 341 107 347 109
rect 341 105 343 107
rect 345 105 347 107
rect 341 103 347 105
rect 342 98 344 103
rect 352 98 354 113
rect 358 112 364 114
rect 358 110 360 112
rect 362 110 364 112
rect 358 108 364 110
rect 359 98 361 108
rect 369 100 371 118
rect 392 100 394 118
rect 402 114 404 128
rect 409 125 411 128
rect 409 123 415 125
rect 409 121 411 123
rect 413 121 415 123
rect 409 119 415 121
rect 419 115 421 128
rect 399 112 405 114
rect 399 110 401 112
rect 403 110 405 112
rect 399 108 405 110
rect 409 113 421 115
rect 426 119 428 128
rect 426 117 432 119
rect 426 115 428 117
rect 430 115 432 117
rect 426 113 432 115
rect 318 95 320 97
rect 322 95 324 97
rect 318 93 324 95
rect 283 84 285 89
rect 293 84 295 89
rect 303 87 305 91
rect 256 78 258 82
rect 402 98 404 108
rect 409 98 411 113
rect 416 107 422 109
rect 416 105 418 107
rect 420 105 422 107
rect 416 103 422 105
rect 419 98 421 103
rect 426 98 428 113
rect 436 110 438 128
rect 503 134 505 144
rect 585 144 610 146
rect 525 131 527 136
rect 459 124 461 127
rect 458 122 464 124
rect 458 120 460 122
rect 462 120 464 122
rect 458 118 464 120
rect 436 99 438 102
rect 459 100 461 118
rect 469 114 471 128
rect 476 125 478 128
rect 476 123 482 125
rect 476 121 478 123
rect 480 121 482 123
rect 476 119 482 121
rect 486 115 488 128
rect 466 112 472 114
rect 466 110 468 112
rect 470 110 472 112
rect 466 108 472 110
rect 476 113 488 115
rect 493 119 495 128
rect 493 117 499 119
rect 493 115 495 117
rect 497 115 499 117
rect 493 113 499 115
rect 436 97 445 99
rect 439 95 441 97
rect 443 95 445 97
rect 439 93 445 95
rect 469 98 471 108
rect 476 98 478 113
rect 483 107 489 109
rect 483 105 485 107
rect 487 105 489 107
rect 483 103 489 105
rect 486 98 488 103
rect 493 98 495 113
rect 503 110 505 128
rect 535 128 537 133
rect 545 128 547 133
rect 568 139 570 144
rect 575 139 577 144
rect 585 136 587 144
rect 595 136 597 140
rect 608 136 610 144
rect 608 134 613 136
rect 611 131 613 134
rect 525 119 527 122
rect 535 119 537 122
rect 525 117 531 119
rect 525 115 527 117
rect 529 115 531 117
rect 525 113 531 115
rect 535 117 541 119
rect 535 115 537 117
rect 539 115 541 117
rect 535 113 541 115
rect 525 110 527 113
rect 503 99 505 102
rect 503 97 512 99
rect 506 95 508 97
rect 510 95 512 97
rect 506 93 512 95
rect 538 103 540 113
rect 545 112 547 122
rect 568 118 570 127
rect 575 124 577 127
rect 575 122 579 124
rect 585 123 587 127
rect 595 124 597 127
rect 577 119 579 122
rect 595 122 604 124
rect 595 120 600 122
rect 602 120 604 122
rect 567 116 573 118
rect 567 114 569 116
rect 571 114 573 116
rect 567 112 573 114
rect 577 117 583 119
rect 577 115 579 117
rect 581 115 583 117
rect 577 113 583 115
rect 595 118 604 120
rect 595 114 597 118
rect 611 114 613 122
rect 545 110 551 112
rect 545 108 547 110
rect 549 108 551 110
rect 567 109 569 112
rect 577 109 579 113
rect 587 112 597 114
rect 603 112 616 114
rect 587 109 589 112
rect 603 109 605 112
rect 614 111 616 112
rect 614 109 620 111
rect 545 106 551 108
rect 545 103 547 106
rect 525 87 527 92
rect 335 78 337 82
rect 342 78 344 82
rect 352 78 354 82
rect 359 78 361 82
rect 369 78 371 82
rect 392 78 394 82
rect 402 78 404 82
rect 409 78 411 82
rect 419 78 421 82
rect 426 78 428 82
rect 459 78 461 82
rect 469 78 471 82
rect 476 78 478 82
rect 486 78 488 82
rect 493 78 495 82
rect 577 87 579 91
rect 587 87 589 91
rect 538 78 540 82
rect 545 78 547 82
rect 567 78 569 82
rect 614 107 616 109
rect 618 107 620 109
rect 614 105 620 107
rect 603 78 605 82
rect 23 70 25 74
rect 30 70 32 74
rect 10 60 12 65
rect 107 70 109 74
rect 59 61 61 65
rect 69 63 71 68
rect 79 63 81 68
rect 10 39 12 42
rect 23 39 25 49
rect 30 46 32 49
rect 30 44 36 46
rect 30 42 32 44
rect 34 42 36 44
rect 30 40 36 42
rect 10 37 16 39
rect 10 35 12 37
rect 14 35 16 37
rect 10 33 16 35
rect 20 37 26 39
rect 20 35 22 37
rect 24 35 26 37
rect 20 33 26 35
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 40
rect 59 39 61 43
rect 69 39 71 50
rect 79 47 81 50
rect 79 45 85 47
rect 79 43 81 45
rect 83 43 85 45
rect 79 41 85 43
rect 92 45 98 47
rect 92 43 94 45
rect 96 43 98 45
rect 143 70 145 74
rect 123 61 125 65
rect 133 61 135 65
rect 221 70 223 74
rect 173 61 175 65
rect 183 63 185 68
rect 193 63 195 68
rect 92 41 98 43
rect 59 37 65 39
rect 59 35 61 37
rect 63 35 65 37
rect 59 33 65 35
rect 69 37 75 39
rect 69 35 71 37
rect 73 35 75 37
rect 69 33 75 35
rect 59 28 61 33
rect 72 28 74 33
rect 79 28 81 41
rect 96 40 98 41
rect 107 40 109 43
rect 123 40 125 43
rect 96 38 109 40
rect 115 38 125 40
rect 133 39 135 43
rect 143 40 145 43
rect 99 30 101 38
rect 115 34 117 38
rect 108 32 117 34
rect 129 37 135 39
rect 129 35 131 37
rect 133 35 135 37
rect 129 33 135 35
rect 139 38 145 40
rect 139 36 141 38
rect 143 36 145 38
rect 139 34 145 36
rect 173 39 175 43
rect 183 39 185 50
rect 193 47 195 50
rect 193 45 199 47
rect 193 43 195 45
rect 197 43 199 45
rect 193 41 199 43
rect 206 45 212 47
rect 206 43 208 45
rect 210 43 212 45
rect 257 70 259 74
rect 237 61 239 65
rect 247 61 249 65
rect 336 70 338 74
rect 343 70 345 74
rect 353 70 355 74
rect 360 70 362 74
rect 370 70 372 74
rect 393 70 395 74
rect 403 70 405 74
rect 410 70 412 74
rect 420 70 422 74
rect 427 70 429 74
rect 460 70 462 74
rect 470 70 472 74
rect 477 70 479 74
rect 487 70 489 74
rect 494 70 496 74
rect 284 63 286 68
rect 294 63 296 68
rect 304 61 306 65
rect 284 47 286 50
rect 280 45 286 47
rect 280 43 282 45
rect 284 43 286 45
rect 206 41 212 43
rect 173 37 179 39
rect 173 35 175 37
rect 177 35 179 37
rect 108 30 110 32
rect 112 30 117 32
rect 10 16 12 21
rect 20 19 22 24
rect 30 19 32 24
rect 59 15 61 19
rect 108 28 117 30
rect 133 30 135 33
rect 115 25 117 28
rect 125 25 127 29
rect 133 28 137 30
rect 135 25 137 28
rect 142 25 144 34
rect 173 33 179 35
rect 183 37 189 39
rect 183 35 185 37
rect 187 35 189 37
rect 183 33 189 35
rect 173 28 175 33
rect 186 28 188 33
rect 193 28 195 41
rect 210 40 212 41
rect 221 40 223 43
rect 237 40 239 43
rect 210 38 223 40
rect 229 38 239 40
rect 247 39 249 43
rect 257 40 259 43
rect 280 41 286 43
rect 213 30 215 38
rect 229 34 231 38
rect 222 32 231 34
rect 243 37 249 39
rect 243 35 245 37
rect 247 35 249 37
rect 243 33 249 35
rect 253 38 259 40
rect 253 36 255 38
rect 257 36 259 38
rect 253 34 259 36
rect 222 30 224 32
rect 226 30 231 32
rect 99 18 101 21
rect 72 12 74 17
rect 79 12 81 17
rect 99 16 104 18
rect 102 8 104 16
rect 115 12 117 16
rect 125 8 127 16
rect 173 15 175 19
rect 222 28 231 30
rect 247 30 249 33
rect 229 25 231 28
rect 239 25 241 29
rect 247 28 251 30
rect 249 25 251 28
rect 256 25 258 34
rect 284 28 286 41
rect 294 39 296 50
rect 319 57 325 59
rect 319 55 321 57
rect 323 55 325 57
rect 319 53 328 55
rect 326 50 328 53
rect 304 39 306 43
rect 290 37 296 39
rect 290 35 292 37
rect 294 35 296 37
rect 290 33 296 35
rect 300 37 306 39
rect 300 35 302 37
rect 304 35 306 37
rect 300 33 306 35
rect 291 28 293 33
rect 304 28 306 33
rect 213 18 215 21
rect 135 8 137 13
rect 142 8 144 13
rect 102 6 127 8
rect 186 12 188 17
rect 193 12 195 17
rect 213 16 218 18
rect 216 8 218 16
rect 229 12 231 16
rect 239 8 241 16
rect 326 24 328 42
rect 336 39 338 54
rect 343 49 345 54
rect 342 47 348 49
rect 342 45 344 47
rect 346 45 348 47
rect 342 43 348 45
rect 353 39 355 54
rect 360 44 362 54
rect 440 57 446 59
rect 440 55 442 57
rect 444 55 446 57
rect 332 37 338 39
rect 332 35 334 37
rect 336 35 338 37
rect 332 33 338 35
rect 336 24 338 33
rect 343 37 355 39
rect 359 42 365 44
rect 359 40 361 42
rect 363 40 365 42
rect 359 38 365 40
rect 343 24 345 37
rect 349 31 355 33
rect 349 29 351 31
rect 353 29 355 31
rect 349 27 355 29
rect 353 24 355 27
rect 360 24 362 38
rect 370 34 372 52
rect 393 34 395 52
rect 403 44 405 54
rect 400 42 406 44
rect 400 40 402 42
rect 404 40 406 42
rect 400 38 406 40
rect 410 39 412 54
rect 420 49 422 54
rect 417 47 423 49
rect 417 45 419 47
rect 421 45 423 47
rect 417 43 423 45
rect 427 39 429 54
rect 437 53 446 55
rect 437 50 439 53
rect 539 70 541 74
rect 546 70 548 74
rect 568 70 570 74
rect 526 60 528 65
rect 507 57 513 59
rect 507 55 509 57
rect 511 55 513 57
rect 367 32 373 34
rect 367 30 369 32
rect 371 30 373 32
rect 367 28 373 30
rect 392 32 398 34
rect 392 30 394 32
rect 396 30 398 32
rect 392 28 398 30
rect 370 25 372 28
rect 393 25 395 28
rect 249 8 251 13
rect 256 8 258 13
rect 284 12 286 17
rect 291 12 293 17
rect 216 6 241 8
rect 304 15 306 19
rect 326 8 328 18
rect 403 24 405 38
rect 410 37 422 39
rect 410 31 416 33
rect 410 29 412 31
rect 414 29 416 31
rect 410 27 416 29
rect 410 24 412 27
rect 420 24 422 37
rect 427 37 433 39
rect 427 35 429 37
rect 431 35 433 37
rect 427 33 433 35
rect 427 24 429 33
rect 437 24 439 42
rect 460 34 462 52
rect 470 44 472 54
rect 467 42 473 44
rect 467 40 469 42
rect 471 40 473 42
rect 467 38 473 40
rect 477 39 479 54
rect 487 49 489 54
rect 484 47 490 49
rect 484 45 486 47
rect 488 45 490 47
rect 484 43 490 45
rect 494 39 496 54
rect 504 53 513 55
rect 504 50 506 53
rect 459 32 465 34
rect 459 30 461 32
rect 463 30 465 32
rect 459 28 465 30
rect 460 25 462 28
rect 336 12 338 16
rect 343 8 345 16
rect 353 11 355 16
rect 360 11 362 16
rect 370 11 372 16
rect 393 11 395 16
rect 403 11 405 16
rect 410 11 412 16
rect 326 6 345 8
rect 420 8 422 16
rect 427 12 429 16
rect 437 8 439 18
rect 470 24 472 38
rect 477 37 489 39
rect 477 31 483 33
rect 477 29 479 31
rect 481 29 483 31
rect 477 27 483 29
rect 477 24 479 27
rect 487 24 489 37
rect 494 37 500 39
rect 494 35 496 37
rect 498 35 500 37
rect 494 33 500 35
rect 494 24 496 33
rect 504 24 506 42
rect 526 39 528 42
rect 539 39 541 49
rect 546 46 548 49
rect 546 44 552 46
rect 546 42 548 44
rect 550 42 552 44
rect 604 70 606 74
rect 578 61 580 65
rect 588 61 590 65
rect 615 45 621 47
rect 615 43 617 45
rect 619 43 621 45
rect 546 40 552 42
rect 568 40 570 43
rect 526 37 532 39
rect 526 35 528 37
rect 530 35 532 37
rect 526 33 532 35
rect 536 37 542 39
rect 536 35 538 37
rect 540 35 542 37
rect 536 33 542 35
rect 526 30 528 33
rect 536 30 538 33
rect 546 30 548 40
rect 568 38 574 40
rect 568 36 570 38
rect 572 36 574 38
rect 568 34 574 36
rect 578 39 580 43
rect 588 40 590 43
rect 604 40 606 43
rect 615 41 621 43
rect 615 40 617 41
rect 578 37 584 39
rect 588 38 598 40
rect 604 38 617 40
rect 578 35 580 37
rect 582 35 584 37
rect 569 25 571 34
rect 578 33 584 35
rect 596 34 598 38
rect 578 30 580 33
rect 576 28 580 30
rect 596 32 605 34
rect 596 30 601 32
rect 603 30 605 32
rect 612 30 614 38
rect 576 25 578 28
rect 586 25 588 29
rect 596 28 605 30
rect 596 25 598 28
rect 460 11 462 16
rect 470 11 472 16
rect 477 11 479 16
rect 420 6 439 8
rect 487 8 489 16
rect 494 12 496 16
rect 504 8 506 18
rect 526 16 528 21
rect 536 19 538 24
rect 546 19 548 24
rect 487 6 506 8
rect 612 18 614 21
rect 609 16 614 18
rect 569 8 571 13
rect 576 8 578 13
rect 586 8 588 16
rect 596 12 598 16
rect 609 8 611 16
rect 586 6 611 8
<< ndif >>
rect 13 139 19 141
rect 13 137 15 139
rect 17 137 19 139
rect 13 135 19 137
rect 32 139 38 141
rect 62 143 69 145
rect 62 141 64 143
rect 66 141 69 143
rect 32 137 34 139
rect 36 137 38 139
rect 32 135 38 137
rect 13 131 17 135
rect 4 128 9 131
rect 2 126 9 128
rect 2 124 4 126
rect 6 124 9 126
rect 2 122 9 124
rect 11 128 17 131
rect 33 128 38 135
rect 62 135 69 141
rect 145 143 151 145
rect 145 141 147 143
rect 149 141 151 143
rect 145 139 151 141
rect 176 143 183 145
rect 176 141 178 143
rect 180 141 183 143
rect 129 136 134 139
rect 62 133 71 135
rect 11 122 19 128
rect 21 126 29 128
rect 21 124 24 126
rect 26 124 29 126
rect 21 122 29 124
rect 31 122 38 128
rect 51 131 58 133
rect 51 129 53 131
rect 55 129 58 131
rect 51 127 58 129
rect 53 124 58 127
rect 60 124 71 133
rect 73 124 78 135
rect 80 133 87 135
rect 80 131 83 133
rect 85 131 87 133
rect 105 134 114 136
rect 105 132 107 134
rect 109 132 114 134
rect 105 131 114 132
rect 80 129 87 131
rect 80 124 85 129
rect 93 128 98 131
rect 91 126 98 128
rect 91 124 93 126
rect 95 124 98 126
rect 91 122 98 124
rect 100 127 114 131
rect 116 131 124 136
rect 116 129 119 131
rect 121 129 124 131
rect 116 127 124 129
rect 126 133 134 136
rect 126 131 129 133
rect 131 131 134 133
rect 126 127 134 131
rect 136 127 141 139
rect 143 127 151 139
rect 176 135 183 141
rect 259 143 265 145
rect 259 141 261 143
rect 263 141 265 143
rect 259 139 265 141
rect 294 143 301 145
rect 294 141 297 143
rect 299 141 301 143
rect 243 136 248 139
rect 176 133 185 135
rect 165 131 172 133
rect 165 129 167 131
rect 169 129 172 131
rect 165 127 172 129
rect 100 122 105 127
rect 167 124 172 127
rect 174 124 185 133
rect 187 124 192 135
rect 194 133 201 135
rect 194 131 197 133
rect 199 131 201 133
rect 219 134 228 136
rect 219 132 221 134
rect 223 132 228 134
rect 219 131 228 132
rect 194 129 201 131
rect 194 124 199 129
rect 207 128 212 131
rect 205 126 212 128
rect 205 124 207 126
rect 209 124 212 126
rect 205 122 212 124
rect 214 127 228 131
rect 230 131 238 136
rect 230 129 233 131
rect 235 129 238 131
rect 230 127 238 129
rect 240 133 248 136
rect 240 131 243 133
rect 245 131 248 133
rect 240 127 248 131
rect 250 127 255 139
rect 257 127 265 139
rect 294 135 301 141
rect 276 133 283 135
rect 276 131 278 133
rect 280 131 283 133
rect 276 129 283 131
rect 214 122 219 127
rect 278 124 283 129
rect 285 124 290 135
rect 292 133 301 135
rect 329 134 335 136
rect 292 124 303 133
rect 305 131 312 133
rect 305 129 308 131
rect 310 129 312 131
rect 305 127 312 129
rect 318 132 325 134
rect 318 130 320 132
rect 322 130 325 132
rect 318 128 325 130
rect 327 132 335 134
rect 327 130 330 132
rect 332 130 335 132
rect 327 128 335 130
rect 337 128 342 136
rect 344 134 352 136
rect 344 132 347 134
rect 349 132 352 134
rect 344 128 352 132
rect 354 128 359 136
rect 361 134 369 136
rect 361 132 364 134
rect 366 132 369 134
rect 361 128 369 132
rect 305 124 310 127
rect 364 127 369 128
rect 371 133 376 136
rect 387 133 392 136
rect 371 131 378 133
rect 371 129 374 131
rect 376 129 378 131
rect 371 127 378 129
rect 385 131 392 133
rect 385 129 387 131
rect 389 129 392 131
rect 385 127 392 129
rect 394 134 402 136
rect 394 132 397 134
rect 399 132 402 134
rect 394 128 402 132
rect 404 128 409 136
rect 411 134 419 136
rect 411 132 414 134
rect 416 132 419 134
rect 411 128 419 132
rect 421 128 426 136
rect 428 134 434 136
rect 428 132 436 134
rect 428 130 431 132
rect 433 130 436 132
rect 428 128 436 130
rect 438 132 445 134
rect 454 133 459 136
rect 438 130 441 132
rect 443 130 445 132
rect 438 128 445 130
rect 452 131 459 133
rect 452 129 454 131
rect 456 129 459 131
rect 394 127 399 128
rect 452 127 459 129
rect 461 134 469 136
rect 461 132 464 134
rect 466 132 469 134
rect 461 128 469 132
rect 471 128 476 136
rect 478 134 486 136
rect 478 132 481 134
rect 483 132 486 134
rect 478 128 486 132
rect 488 128 493 136
rect 495 134 501 136
rect 560 143 566 145
rect 560 141 562 143
rect 564 141 566 143
rect 529 139 535 141
rect 529 137 531 139
rect 533 137 535 139
rect 495 132 503 134
rect 495 130 498 132
rect 500 130 503 132
rect 495 128 503 130
rect 505 132 512 134
rect 505 130 508 132
rect 510 130 512 132
rect 529 135 535 137
rect 548 139 554 141
rect 548 137 550 139
rect 552 137 554 139
rect 548 135 554 137
rect 529 131 533 135
rect 505 128 512 130
rect 520 128 525 131
rect 461 127 466 128
rect 518 126 525 128
rect 518 124 520 126
rect 522 124 525 126
rect 518 122 525 124
rect 527 128 533 131
rect 549 128 554 135
rect 527 122 535 128
rect 537 126 545 128
rect 537 124 540 126
rect 542 124 545 126
rect 537 122 545 124
rect 547 122 554 128
rect 560 139 566 141
rect 560 127 568 139
rect 570 127 575 139
rect 577 136 582 139
rect 577 133 585 136
rect 577 131 580 133
rect 582 131 585 133
rect 577 127 585 131
rect 587 131 595 136
rect 587 129 590 131
rect 592 129 595 131
rect 587 127 595 129
rect 597 134 606 136
rect 597 132 602 134
rect 604 132 606 134
rect 597 131 606 132
rect 597 127 611 131
rect 606 122 611 127
rect 613 128 618 131
rect 613 126 620 128
rect 613 124 616 126
rect 618 124 620 126
rect 613 122 620 124
rect 3 28 10 30
rect 3 26 5 28
rect 7 26 10 28
rect 3 24 10 26
rect 5 21 10 24
rect 12 24 20 30
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 24 30 26
rect 32 24 39 30
rect 92 28 99 30
rect 54 25 59 28
rect 12 21 18 24
rect 14 17 18 21
rect 34 17 39 24
rect 52 23 59 25
rect 52 21 54 23
rect 56 21 59 23
rect 52 19 59 21
rect 61 19 72 28
rect 14 15 20 17
rect 14 13 16 15
rect 18 13 20 15
rect 14 11 20 13
rect 33 15 39 17
rect 63 17 72 19
rect 74 17 79 28
rect 81 23 86 28
rect 92 26 94 28
rect 96 26 99 28
rect 92 24 99 26
rect 81 21 88 23
rect 94 21 99 24
rect 101 25 106 30
rect 206 28 213 30
rect 168 25 173 28
rect 101 21 115 25
rect 81 19 84 21
rect 86 19 88 21
rect 81 17 88 19
rect 106 20 115 21
rect 106 18 108 20
rect 110 18 115 20
rect 33 13 35 15
rect 37 13 39 15
rect 33 11 39 13
rect 63 11 70 17
rect 106 16 115 18
rect 117 23 125 25
rect 117 21 120 23
rect 122 21 125 23
rect 117 16 125 21
rect 127 21 135 25
rect 127 19 130 21
rect 132 19 135 21
rect 127 16 135 19
rect 63 9 65 11
rect 67 9 70 11
rect 63 7 70 9
rect 130 13 135 16
rect 137 13 142 25
rect 144 13 152 25
rect 166 23 173 25
rect 166 21 168 23
rect 170 21 173 23
rect 166 19 173 21
rect 175 19 186 28
rect 177 17 186 19
rect 188 17 193 28
rect 195 23 200 28
rect 206 26 208 28
rect 210 26 213 28
rect 206 24 213 26
rect 195 21 202 23
rect 208 21 213 24
rect 215 25 220 30
rect 215 21 229 25
rect 195 19 198 21
rect 200 19 202 21
rect 195 17 202 19
rect 220 20 229 21
rect 220 18 222 20
rect 224 18 229 20
rect 146 11 152 13
rect 146 9 148 11
rect 150 9 152 11
rect 146 7 152 9
rect 177 11 184 17
rect 220 16 229 18
rect 231 23 239 25
rect 231 21 234 23
rect 236 21 239 23
rect 231 16 239 21
rect 241 21 249 25
rect 241 19 244 21
rect 246 19 249 21
rect 241 16 249 19
rect 177 9 179 11
rect 181 9 184 11
rect 177 7 184 9
rect 244 13 249 16
rect 251 13 256 25
rect 258 13 266 25
rect 279 23 284 28
rect 277 21 284 23
rect 277 19 279 21
rect 281 19 284 21
rect 277 17 284 19
rect 286 17 291 28
rect 293 19 304 28
rect 306 25 311 28
rect 306 23 313 25
rect 365 24 370 25
rect 306 21 309 23
rect 311 21 313 23
rect 306 19 313 21
rect 319 22 326 24
rect 319 20 321 22
rect 323 20 326 22
rect 293 17 302 19
rect 260 11 266 13
rect 260 9 262 11
rect 264 9 266 11
rect 260 7 266 9
rect 295 11 302 17
rect 319 18 326 20
rect 328 22 336 24
rect 328 20 331 22
rect 333 20 336 22
rect 328 18 336 20
rect 295 9 298 11
rect 300 9 302 11
rect 295 7 302 9
rect 330 16 336 18
rect 338 16 343 24
rect 345 20 353 24
rect 345 18 348 20
rect 350 18 353 20
rect 345 16 353 18
rect 355 16 360 24
rect 362 20 370 24
rect 362 18 365 20
rect 367 18 370 20
rect 362 16 370 18
rect 372 23 379 25
rect 372 21 375 23
rect 377 21 379 23
rect 372 19 379 21
rect 386 23 393 25
rect 386 21 388 23
rect 390 21 393 23
rect 386 19 393 21
rect 372 16 377 19
rect 388 16 393 19
rect 395 24 400 25
rect 395 20 403 24
rect 395 18 398 20
rect 400 18 403 20
rect 395 16 403 18
rect 405 16 410 24
rect 412 20 420 24
rect 412 18 415 20
rect 417 18 420 20
rect 412 16 420 18
rect 422 16 427 24
rect 429 22 437 24
rect 429 20 432 22
rect 434 20 437 22
rect 429 18 437 20
rect 439 22 446 24
rect 439 20 442 22
rect 444 20 446 22
rect 439 18 446 20
rect 453 23 460 25
rect 453 21 455 23
rect 457 21 460 23
rect 453 19 460 21
rect 429 16 435 18
rect 455 16 460 19
rect 462 24 467 25
rect 519 28 526 30
rect 519 26 521 28
rect 523 26 526 28
rect 519 24 526 26
rect 462 20 470 24
rect 462 18 465 20
rect 467 18 470 20
rect 462 16 470 18
rect 472 16 477 24
rect 479 20 487 24
rect 479 18 482 20
rect 484 18 487 20
rect 479 16 487 18
rect 489 16 494 24
rect 496 22 504 24
rect 496 20 499 22
rect 501 20 504 22
rect 496 18 504 20
rect 506 22 513 24
rect 506 20 509 22
rect 511 20 513 22
rect 521 21 526 24
rect 528 24 536 30
rect 538 28 546 30
rect 538 26 541 28
rect 543 26 546 28
rect 538 24 546 26
rect 548 24 555 30
rect 607 25 612 30
rect 528 21 534 24
rect 506 18 513 20
rect 496 16 502 18
rect 530 17 534 21
rect 550 17 555 24
rect 530 15 536 17
rect 530 13 532 15
rect 534 13 536 15
rect 530 11 536 13
rect 549 15 555 17
rect 549 13 551 15
rect 553 13 555 15
rect 549 11 555 13
rect 561 13 569 25
rect 571 13 576 25
rect 578 21 586 25
rect 578 19 581 21
rect 583 19 586 21
rect 578 16 586 19
rect 588 23 596 25
rect 588 21 591 23
rect 593 21 596 23
rect 588 16 596 21
rect 598 21 612 25
rect 614 28 621 30
rect 614 26 617 28
rect 619 26 621 28
rect 614 24 621 26
rect 614 21 619 24
rect 598 20 607 21
rect 598 18 603 20
rect 605 18 607 20
rect 598 16 607 18
rect 578 13 583 16
rect 561 11 567 13
rect 561 9 563 11
rect 565 9 567 11
rect 561 7 567 9
<< pdif >>
rect 4 105 9 110
rect 2 103 9 105
rect 2 101 4 103
rect 6 101 9 103
rect 2 96 9 101
rect 2 94 4 96
rect 6 94 9 96
rect 2 92 9 94
rect 11 103 19 110
rect 51 107 58 109
rect 51 105 53 107
rect 55 105 58 107
rect 11 92 22 103
rect 13 86 22 92
rect 13 84 15 86
rect 17 84 22 86
rect 13 82 22 84
rect 24 82 29 103
rect 31 95 36 103
rect 51 100 58 105
rect 51 98 53 100
rect 55 98 58 100
rect 51 96 58 98
rect 31 93 38 95
rect 31 91 34 93
rect 36 91 38 93
rect 53 91 58 96
rect 60 102 66 109
rect 99 107 106 109
rect 99 105 101 107
rect 103 105 106 107
rect 99 103 106 105
rect 60 95 68 102
rect 60 93 63 95
rect 65 93 68 95
rect 60 91 68 93
rect 31 89 38 91
rect 31 82 36 89
rect 62 89 68 91
rect 70 100 78 102
rect 70 98 73 100
rect 75 98 78 100
rect 70 93 78 98
rect 70 91 73 93
rect 75 91 78 93
rect 70 89 78 91
rect 80 93 87 102
rect 80 91 83 93
rect 85 91 87 93
rect 80 89 87 91
rect 101 82 106 103
rect 108 93 122 109
rect 108 91 111 93
rect 113 91 122 93
rect 124 107 132 109
rect 124 105 127 107
rect 129 105 132 107
rect 124 100 132 105
rect 124 98 127 100
rect 129 98 132 100
rect 124 91 132 98
rect 134 100 142 109
rect 134 98 137 100
rect 139 98 142 100
rect 134 91 142 98
rect 108 86 120 91
rect 108 84 111 86
rect 113 84 120 86
rect 108 82 120 84
rect 137 82 142 91
rect 144 94 149 109
rect 165 107 172 109
rect 165 105 167 107
rect 169 105 172 107
rect 165 100 172 105
rect 165 98 167 100
rect 169 98 172 100
rect 165 96 172 98
rect 144 92 151 94
rect 144 90 147 92
rect 149 90 151 92
rect 167 91 172 96
rect 174 102 180 109
rect 213 107 220 109
rect 213 105 215 107
rect 217 105 220 107
rect 213 103 220 105
rect 174 95 182 102
rect 174 93 177 95
rect 179 93 182 95
rect 174 91 182 93
rect 144 88 151 90
rect 144 82 149 88
rect 176 89 182 91
rect 184 100 192 102
rect 184 98 187 100
rect 189 98 192 100
rect 184 93 192 98
rect 184 91 187 93
rect 189 91 192 93
rect 184 89 192 91
rect 194 93 201 102
rect 194 91 197 93
rect 199 91 201 93
rect 194 89 201 91
rect 215 82 220 103
rect 222 93 236 109
rect 222 91 225 93
rect 227 91 236 93
rect 238 107 246 109
rect 238 105 241 107
rect 243 105 246 107
rect 238 100 246 105
rect 238 98 241 100
rect 243 98 246 100
rect 238 91 246 98
rect 248 100 256 109
rect 248 98 251 100
rect 253 98 256 100
rect 248 91 256 98
rect 222 86 234 91
rect 222 84 225 86
rect 227 84 234 86
rect 222 82 234 84
rect 251 82 256 91
rect 258 94 263 109
rect 297 102 303 109
rect 258 92 265 94
rect 258 90 261 92
rect 263 90 265 92
rect 258 88 265 90
rect 276 93 283 102
rect 276 91 278 93
rect 280 91 283 93
rect 276 89 283 91
rect 285 100 293 102
rect 285 98 288 100
rect 290 98 293 100
rect 285 93 293 98
rect 285 91 288 93
rect 290 91 293 93
rect 285 89 293 91
rect 295 95 303 102
rect 295 93 298 95
rect 300 93 303 95
rect 295 91 303 93
rect 305 107 312 109
rect 305 105 308 107
rect 310 105 312 107
rect 305 100 312 105
rect 318 108 325 110
rect 318 106 320 108
rect 322 106 325 108
rect 318 104 325 106
rect 320 102 325 104
rect 327 102 333 110
rect 305 98 308 100
rect 310 98 312 100
rect 305 96 312 98
rect 329 98 333 102
rect 364 98 369 100
rect 305 91 310 96
rect 329 94 335 98
rect 295 89 301 91
rect 258 82 263 88
rect 328 86 335 94
rect 328 84 330 86
rect 332 84 335 86
rect 328 82 335 84
rect 337 82 342 98
rect 344 96 352 98
rect 344 94 347 96
rect 349 94 352 96
rect 344 82 352 94
rect 354 82 359 98
rect 361 86 369 98
rect 361 84 364 86
rect 366 84 369 86
rect 361 82 369 84
rect 371 95 376 100
rect 387 95 392 100
rect 371 93 378 95
rect 371 91 374 93
rect 376 91 378 93
rect 371 89 378 91
rect 385 93 392 95
rect 385 91 387 93
rect 389 91 392 93
rect 385 89 392 91
rect 371 82 376 89
rect 387 82 392 89
rect 394 98 399 100
rect 430 102 436 110
rect 438 108 445 110
rect 438 106 441 108
rect 443 106 445 108
rect 438 104 445 106
rect 438 102 443 104
rect 430 98 434 102
rect 394 86 402 98
rect 394 84 397 86
rect 399 84 402 86
rect 394 82 402 84
rect 404 82 409 98
rect 411 96 419 98
rect 411 94 414 96
rect 416 94 419 96
rect 411 82 419 94
rect 421 82 426 98
rect 428 94 434 98
rect 454 95 459 100
rect 428 86 435 94
rect 452 93 459 95
rect 452 91 454 93
rect 456 91 459 93
rect 452 89 459 91
rect 428 84 431 86
rect 433 84 435 86
rect 428 82 435 84
rect 454 82 459 89
rect 461 98 466 100
rect 497 102 503 110
rect 505 108 512 110
rect 505 106 508 108
rect 510 106 512 108
rect 505 104 512 106
rect 520 105 525 110
rect 505 102 510 104
rect 518 103 525 105
rect 497 98 501 102
rect 461 86 469 98
rect 461 84 464 86
rect 466 84 469 86
rect 461 82 469 84
rect 471 82 476 98
rect 478 96 486 98
rect 478 94 481 96
rect 483 94 486 96
rect 478 82 486 94
rect 488 82 493 98
rect 495 94 501 98
rect 518 101 520 103
rect 522 101 525 103
rect 495 86 502 94
rect 518 96 525 101
rect 518 94 520 96
rect 522 94 525 96
rect 518 92 525 94
rect 527 103 535 110
rect 527 92 538 103
rect 495 84 498 86
rect 500 84 502 86
rect 529 86 538 92
rect 495 82 502 84
rect 529 84 531 86
rect 533 84 538 86
rect 529 82 538 84
rect 540 82 545 103
rect 547 95 552 103
rect 547 93 554 95
rect 562 94 567 109
rect 547 91 550 93
rect 552 91 554 93
rect 547 89 554 91
rect 560 92 567 94
rect 560 90 562 92
rect 564 90 567 92
rect 547 82 552 89
rect 560 88 567 90
rect 562 82 567 88
rect 569 100 577 109
rect 569 98 572 100
rect 574 98 577 100
rect 569 91 577 98
rect 579 107 587 109
rect 579 105 582 107
rect 584 105 587 107
rect 579 100 587 105
rect 579 98 582 100
rect 584 98 587 100
rect 579 91 587 98
rect 589 93 603 109
rect 589 91 598 93
rect 600 91 603 93
rect 569 82 574 91
rect 591 86 603 91
rect 591 84 598 86
rect 600 84 603 86
rect 591 82 603 84
rect 605 107 612 109
rect 605 105 608 107
rect 610 105 612 107
rect 605 103 612 105
rect 605 82 610 103
rect 14 68 23 70
rect 14 66 16 68
rect 18 66 23 68
rect 14 60 23 66
rect 3 58 10 60
rect 3 56 5 58
rect 7 56 10 58
rect 3 51 10 56
rect 3 49 5 51
rect 7 49 10 51
rect 3 47 10 49
rect 5 42 10 47
rect 12 49 23 60
rect 25 49 30 70
rect 32 63 37 70
rect 32 61 39 63
rect 63 61 69 63
rect 32 59 35 61
rect 37 59 39 61
rect 32 57 39 59
rect 32 49 37 57
rect 54 56 59 61
rect 52 54 59 56
rect 52 52 54 54
rect 56 52 59 54
rect 12 42 20 49
rect 52 47 59 52
rect 52 45 54 47
rect 56 45 59 47
rect 52 43 59 45
rect 61 59 69 61
rect 61 57 64 59
rect 66 57 69 59
rect 61 50 69 57
rect 71 61 79 63
rect 71 59 74 61
rect 76 59 79 61
rect 71 54 79 59
rect 71 52 74 54
rect 76 52 79 54
rect 71 50 79 52
rect 81 61 88 63
rect 81 59 84 61
rect 86 59 88 61
rect 81 50 88 59
rect 61 43 67 50
rect 102 49 107 70
rect 100 47 107 49
rect 100 45 102 47
rect 104 45 107 47
rect 100 43 107 45
rect 109 68 121 70
rect 109 66 112 68
rect 114 66 121 68
rect 109 61 121 66
rect 138 61 143 70
rect 109 59 112 61
rect 114 59 123 61
rect 109 43 123 59
rect 125 54 133 61
rect 125 52 128 54
rect 130 52 133 54
rect 125 47 133 52
rect 125 45 128 47
rect 130 45 133 47
rect 125 43 133 45
rect 135 54 143 61
rect 135 52 138 54
rect 140 52 143 54
rect 135 43 143 52
rect 145 64 150 70
rect 145 62 152 64
rect 145 60 148 62
rect 150 60 152 62
rect 177 61 183 63
rect 145 58 152 60
rect 145 43 150 58
rect 168 56 173 61
rect 166 54 173 56
rect 166 52 168 54
rect 170 52 173 54
rect 166 47 173 52
rect 166 45 168 47
rect 170 45 173 47
rect 166 43 173 45
rect 175 59 183 61
rect 175 57 178 59
rect 180 57 183 59
rect 175 50 183 57
rect 185 61 193 63
rect 185 59 188 61
rect 190 59 193 61
rect 185 54 193 59
rect 185 52 188 54
rect 190 52 193 54
rect 185 50 193 52
rect 195 61 202 63
rect 195 59 198 61
rect 200 59 202 61
rect 195 50 202 59
rect 175 43 181 50
rect 216 49 221 70
rect 214 47 221 49
rect 214 45 216 47
rect 218 45 221 47
rect 214 43 221 45
rect 223 68 235 70
rect 223 66 226 68
rect 228 66 235 68
rect 223 61 235 66
rect 252 61 257 70
rect 223 59 226 61
rect 228 59 237 61
rect 223 43 237 59
rect 239 54 247 61
rect 239 52 242 54
rect 244 52 247 54
rect 239 47 247 52
rect 239 45 242 47
rect 244 45 247 47
rect 239 43 247 45
rect 249 54 257 61
rect 249 52 252 54
rect 254 52 257 54
rect 249 43 257 52
rect 259 64 264 70
rect 259 62 266 64
rect 329 68 336 70
rect 329 66 331 68
rect 333 66 336 68
rect 259 60 262 62
rect 264 60 266 62
rect 259 58 266 60
rect 277 61 284 63
rect 277 59 279 61
rect 281 59 284 61
rect 259 43 264 58
rect 277 50 284 59
rect 286 61 294 63
rect 286 59 289 61
rect 291 59 294 61
rect 286 54 294 59
rect 286 52 289 54
rect 291 52 294 54
rect 286 50 294 52
rect 296 61 302 63
rect 296 59 304 61
rect 296 57 299 59
rect 301 57 304 59
rect 296 50 304 57
rect 298 43 304 50
rect 306 56 311 61
rect 329 58 336 66
rect 306 54 313 56
rect 306 52 309 54
rect 311 52 313 54
rect 306 47 313 52
rect 330 54 336 58
rect 338 54 343 70
rect 345 58 353 70
rect 345 56 348 58
rect 350 56 353 58
rect 345 54 353 56
rect 355 54 360 70
rect 362 68 370 70
rect 362 66 365 68
rect 367 66 370 68
rect 362 54 370 66
rect 330 50 334 54
rect 321 48 326 50
rect 306 45 309 47
rect 311 45 313 47
rect 306 43 313 45
rect 319 46 326 48
rect 319 44 321 46
rect 323 44 326 46
rect 319 42 326 44
rect 328 42 334 50
rect 365 52 370 54
rect 372 63 377 70
rect 388 63 393 70
rect 372 61 379 63
rect 372 59 375 61
rect 377 59 379 61
rect 372 57 379 59
rect 386 61 393 63
rect 386 59 388 61
rect 390 59 393 61
rect 386 57 393 59
rect 372 52 377 57
rect 388 52 393 57
rect 395 68 403 70
rect 395 66 398 68
rect 400 66 403 68
rect 395 54 403 66
rect 405 54 410 70
rect 412 58 420 70
rect 412 56 415 58
rect 417 56 420 58
rect 412 54 420 56
rect 422 54 427 70
rect 429 68 436 70
rect 429 66 432 68
rect 434 66 436 68
rect 429 58 436 66
rect 455 63 460 70
rect 453 61 460 63
rect 453 59 455 61
rect 457 59 460 61
rect 429 54 435 58
rect 453 57 460 59
rect 395 52 400 54
rect 431 50 435 54
rect 455 52 460 57
rect 462 68 470 70
rect 462 66 465 68
rect 467 66 470 68
rect 462 54 470 66
rect 472 54 477 70
rect 479 58 487 70
rect 479 56 482 58
rect 484 56 487 58
rect 479 54 487 56
rect 489 54 494 70
rect 496 68 503 70
rect 496 66 499 68
rect 501 66 503 68
rect 530 68 539 70
rect 496 58 503 66
rect 530 66 532 68
rect 534 66 539 68
rect 530 60 539 66
rect 496 54 502 58
rect 462 52 467 54
rect 431 42 437 50
rect 439 48 444 50
rect 439 46 446 48
rect 439 44 442 46
rect 444 44 446 46
rect 439 42 446 44
rect 498 50 502 54
rect 519 58 526 60
rect 519 56 521 58
rect 523 56 526 58
rect 519 51 526 56
rect 498 42 504 50
rect 506 48 511 50
rect 519 49 521 51
rect 523 49 526 51
rect 506 46 513 48
rect 519 47 526 49
rect 506 44 509 46
rect 511 44 513 46
rect 506 42 513 44
rect 521 42 526 47
rect 528 49 539 60
rect 541 49 546 70
rect 548 63 553 70
rect 563 64 568 70
rect 548 61 555 63
rect 548 59 551 61
rect 553 59 555 61
rect 548 57 555 59
rect 561 62 568 64
rect 561 60 563 62
rect 565 60 568 62
rect 561 58 568 60
rect 548 49 553 57
rect 528 42 536 49
rect 563 43 568 58
rect 570 61 575 70
rect 592 68 604 70
rect 592 66 599 68
rect 601 66 604 68
rect 592 61 604 66
rect 570 54 578 61
rect 570 52 573 54
rect 575 52 578 54
rect 570 43 578 52
rect 580 54 588 61
rect 580 52 583 54
rect 585 52 588 54
rect 580 47 588 52
rect 580 45 583 47
rect 585 45 588 47
rect 580 43 588 45
rect 590 59 599 61
rect 601 59 604 61
rect 590 43 604 59
rect 606 49 611 70
rect 606 47 613 49
rect 606 45 609 47
rect 611 45 613 47
rect 606 43 613 45
<< alu1 >>
rect -2 143 628 148
rect -2 141 5 143
rect 7 141 54 143
rect 56 141 64 143
rect 66 141 94 143
rect 96 141 147 143
rect 149 141 168 143
rect 170 141 178 143
rect 180 141 208 143
rect 210 141 261 143
rect 263 141 297 143
rect 299 141 307 143
rect 309 141 521 143
rect 523 141 562 143
rect 564 141 615 143
rect 617 141 628 143
rect -2 140 628 141
rect 51 131 63 135
rect 51 129 53 131
rect 55 129 63 131
rect 127 133 151 134
rect 2 126 7 128
rect 2 124 4 126
rect 6 124 7 126
rect 2 122 7 124
rect 2 103 6 122
rect 34 118 38 127
rect 2 101 4 103
rect 2 96 6 101
rect 2 94 4 96
rect 17 117 38 118
rect 17 115 21 117
rect 23 115 35 117
rect 37 115 38 117
rect 17 114 38 115
rect 17 108 31 110
rect 33 108 38 110
rect 17 106 38 108
rect 34 104 38 106
rect 51 109 55 129
rect 127 131 129 133
rect 131 131 151 133
rect 127 130 151 131
rect 75 126 80 127
rect 75 124 76 126
rect 78 124 80 126
rect 75 118 80 124
rect 51 107 56 109
rect 51 105 53 107
rect 55 105 56 107
rect 51 104 56 105
rect 34 100 56 104
rect 34 97 38 100
rect 51 98 53 100
rect 55 98 56 100
rect 66 117 80 118
rect 66 115 70 117
rect 72 115 80 117
rect 66 114 80 115
rect 99 126 112 127
rect 99 124 101 126
rect 103 124 112 126
rect 99 122 112 124
rect 99 121 109 122
rect 107 120 109 121
rect 111 120 112 122
rect 74 109 87 110
rect 74 107 80 109
rect 82 107 87 109
rect 74 106 87 107
rect 51 96 56 98
rect 2 90 15 94
rect 2 89 6 90
rect 83 102 87 106
rect 83 100 84 102
rect 86 100 87 102
rect 83 97 87 100
rect 91 109 96 111
rect 91 107 93 109
rect 95 107 96 109
rect 91 102 96 107
rect 107 113 112 120
rect 147 125 151 130
rect 147 123 148 125
rect 150 123 151 125
rect 91 100 93 102
rect 95 100 96 102
rect 91 95 96 100
rect 91 89 103 95
rect 147 102 151 123
rect 135 100 151 102
rect 135 98 137 100
rect 139 98 151 100
rect 135 97 151 98
rect 165 131 177 135
rect 165 129 167 131
rect 169 129 177 131
rect 241 133 265 134
rect 165 117 169 129
rect 241 131 243 133
rect 245 131 265 133
rect 241 130 265 131
rect 165 115 166 117
rect 168 115 169 117
rect 165 109 169 115
rect 189 126 194 127
rect 189 124 190 126
rect 192 124 194 126
rect 189 118 194 124
rect 165 107 170 109
rect 165 105 167 107
rect 169 105 170 107
rect 165 100 170 105
rect 165 98 167 100
rect 169 98 170 100
rect 180 117 194 118
rect 180 115 184 117
rect 186 115 194 117
rect 180 114 194 115
rect 213 126 226 127
rect 213 124 215 126
rect 217 124 226 126
rect 213 122 226 124
rect 213 121 223 122
rect 221 120 223 121
rect 225 120 226 122
rect 188 109 201 110
rect 188 107 194 109
rect 196 107 201 109
rect 188 106 201 107
rect 165 96 170 98
rect 197 102 201 106
rect 197 100 198 102
rect 200 100 201 102
rect 197 97 201 100
rect 205 109 210 111
rect 205 107 207 109
rect 209 107 210 109
rect 205 102 210 107
rect 221 113 226 120
rect 205 100 207 102
rect 209 100 210 102
rect 205 95 210 100
rect 205 89 217 95
rect 261 110 265 130
rect 283 118 288 127
rect 300 131 312 135
rect 300 129 308 131
rect 310 129 312 131
rect 283 117 297 118
rect 283 115 291 117
rect 293 115 297 117
rect 283 114 297 115
rect 261 108 262 110
rect 264 108 265 110
rect 261 102 265 108
rect 249 100 265 102
rect 249 98 251 100
rect 253 98 265 100
rect 249 97 265 98
rect 276 109 289 110
rect 276 107 281 109
rect 283 107 289 109
rect 276 106 289 107
rect 276 97 280 106
rect 308 125 312 129
rect 308 123 309 125
rect 311 123 312 125
rect 308 109 312 123
rect 307 107 312 109
rect 307 105 308 107
rect 310 105 312 107
rect 374 133 378 135
rect 373 131 378 133
rect 373 129 374 131
rect 376 129 378 131
rect 373 127 378 129
rect 325 125 338 126
rect 325 123 326 125
rect 328 123 338 125
rect 325 122 338 123
rect 332 117 338 122
rect 332 115 333 117
rect 335 115 338 117
rect 332 113 338 115
rect 358 112 362 119
rect 358 111 360 112
rect 350 110 360 111
rect 350 109 362 110
rect 350 107 351 109
rect 353 107 362 109
rect 350 105 362 107
rect 307 100 312 105
rect 307 98 308 100
rect 310 98 312 100
rect 307 96 312 98
rect 318 101 331 102
rect 318 99 328 101
rect 330 99 331 101
rect 318 98 331 99
rect 318 97 323 98
rect 374 117 378 127
rect 374 115 375 117
rect 377 115 378 117
rect 318 95 320 97
rect 322 95 323 97
rect 318 89 323 95
rect 374 94 378 115
rect 365 93 378 94
rect 365 91 374 93
rect 376 91 378 93
rect 365 90 378 91
rect 385 133 389 135
rect 385 131 390 133
rect 385 129 387 131
rect 389 129 390 131
rect 452 133 456 135
rect 385 127 390 129
rect 385 94 389 127
rect 425 125 438 126
rect 401 117 405 119
rect 401 115 402 117
rect 404 115 405 117
rect 401 112 405 115
rect 403 111 405 112
rect 403 110 413 111
rect 401 105 413 110
rect 425 123 433 125
rect 435 123 438 125
rect 425 122 438 123
rect 425 117 431 122
rect 425 115 428 117
rect 430 115 431 117
rect 425 113 431 115
rect 452 131 457 133
rect 452 129 454 131
rect 456 129 457 131
rect 560 133 584 134
rect 452 127 457 129
rect 452 125 456 127
rect 452 123 453 125
rect 455 123 456 125
rect 492 125 505 126
rect 432 98 445 102
rect 440 97 445 98
rect 385 93 398 94
rect 440 95 441 97
rect 443 95 445 97
rect 385 91 387 93
rect 389 91 398 93
rect 385 90 398 91
rect 440 89 445 95
rect 452 94 456 123
rect 468 112 472 119
rect 470 111 472 112
rect 470 110 480 111
rect 468 108 476 110
rect 478 108 480 110
rect 468 105 480 108
rect 492 123 501 125
rect 503 123 505 125
rect 492 122 505 123
rect 492 117 498 122
rect 492 115 495 117
rect 497 115 498 117
rect 492 113 498 115
rect 560 131 580 133
rect 582 131 584 133
rect 560 130 584 131
rect 518 126 523 128
rect 518 124 520 126
rect 522 124 523 126
rect 518 122 523 124
rect 518 109 522 122
rect 518 107 519 109
rect 521 107 522 109
rect 518 103 522 107
rect 550 118 554 127
rect 499 101 512 102
rect 499 99 500 101
rect 502 99 512 101
rect 499 98 512 99
rect 507 97 512 98
rect 452 93 465 94
rect 507 95 508 97
rect 510 95 512 97
rect 452 91 454 93
rect 456 91 465 93
rect 452 90 465 91
rect 507 89 512 95
rect 518 101 520 103
rect 518 96 522 101
rect 518 94 520 96
rect 533 117 554 118
rect 533 115 537 117
rect 539 115 554 117
rect 533 114 554 115
rect 560 125 564 130
rect 560 123 561 125
rect 563 123 564 125
rect 533 108 547 110
rect 549 108 554 110
rect 533 106 554 108
rect 550 97 554 106
rect 560 102 564 123
rect 599 122 612 127
rect 599 120 600 122
rect 602 121 612 122
rect 602 120 604 121
rect 560 100 576 102
rect 560 98 572 100
rect 574 98 576 100
rect 560 97 576 98
rect 599 113 604 120
rect 615 109 620 111
rect 615 107 616 109
rect 618 107 620 109
rect 518 90 531 94
rect 615 95 620 107
rect 518 89 522 90
rect 608 89 620 95
rect -2 83 628 84
rect -2 81 5 83
rect 7 81 54 83
rect 56 81 127 83
rect 129 81 168 83
rect 170 81 241 83
rect 243 81 307 83
rect 309 81 521 83
rect 523 81 582 83
rect 584 81 628 83
rect -2 76 628 81
rect -1 71 629 76
rect -1 69 6 71
rect 8 69 55 71
rect 57 69 128 71
rect 130 69 169 71
rect 171 69 242 71
rect 244 69 308 71
rect 310 69 522 71
rect 524 69 583 71
rect 585 69 629 71
rect -1 68 629 69
rect 3 62 7 63
rect 3 58 16 62
rect 3 56 5 58
rect 3 51 7 56
rect 3 49 5 51
rect 3 46 7 49
rect 35 52 39 55
rect 52 54 57 56
rect 52 52 54 54
rect 56 52 57 54
rect 92 57 104 63
rect 3 44 4 46
rect 6 44 7 46
rect 3 30 7 44
rect 35 48 57 52
rect 35 46 39 48
rect 18 44 39 46
rect 18 42 32 44
rect 34 42 39 44
rect 52 47 57 48
rect 52 45 54 47
rect 56 45 57 47
rect 52 43 57 45
rect 84 52 88 55
rect 84 50 85 52
rect 87 50 88 52
rect 3 28 8 30
rect 3 26 5 28
rect 7 26 8 28
rect 3 24 8 26
rect 18 37 39 38
rect 18 35 22 37
rect 24 35 36 37
rect 38 35 39 37
rect 18 34 39 35
rect 35 25 39 34
rect 52 23 56 43
rect 84 46 88 50
rect 75 45 88 46
rect 75 43 81 45
rect 83 43 88 45
rect 75 42 88 43
rect 92 52 97 57
rect 92 50 94 52
rect 96 50 97 52
rect 92 45 97 50
rect 92 43 94 45
rect 96 43 97 45
rect 92 41 97 43
rect 67 37 81 38
rect 67 35 71 37
rect 73 35 81 37
rect 67 34 81 35
rect 52 21 54 23
rect 56 21 64 23
rect 52 17 64 21
rect 76 28 81 34
rect 76 26 77 28
rect 79 26 81 28
rect 76 25 81 26
rect 108 32 113 39
rect 136 54 152 55
rect 136 52 138 54
rect 140 52 152 54
rect 136 50 152 52
rect 108 31 110 32
rect 100 30 110 31
rect 112 30 113 32
rect 100 28 113 30
rect 100 26 102 28
rect 104 26 113 28
rect 100 25 113 26
rect 148 29 152 50
rect 148 27 149 29
rect 151 27 152 29
rect 148 22 152 27
rect 128 21 152 22
rect 128 19 130 21
rect 132 19 152 21
rect 128 18 152 19
rect 166 54 171 56
rect 166 52 168 54
rect 170 52 171 54
rect 206 57 218 63
rect 166 47 171 52
rect 166 45 168 47
rect 170 45 171 47
rect 166 43 171 45
rect 198 52 202 55
rect 198 50 199 52
rect 201 50 202 52
rect 166 37 170 43
rect 166 35 167 37
rect 169 35 170 37
rect 166 23 170 35
rect 198 46 202 50
rect 189 45 202 46
rect 189 43 195 45
rect 197 43 202 45
rect 189 42 202 43
rect 206 52 211 57
rect 206 50 208 52
rect 210 50 211 52
rect 206 45 211 50
rect 206 43 208 45
rect 210 43 211 45
rect 206 41 211 43
rect 181 37 195 38
rect 181 35 185 37
rect 187 35 195 37
rect 181 34 195 35
rect 166 21 168 23
rect 170 21 178 23
rect 166 17 178 21
rect 190 28 195 34
rect 190 26 191 28
rect 193 26 195 28
rect 190 25 195 26
rect 222 32 227 39
rect 250 54 266 55
rect 250 52 252 54
rect 254 52 266 54
rect 250 50 266 52
rect 262 44 266 50
rect 262 42 263 44
rect 265 42 266 44
rect 277 46 281 55
rect 319 57 324 63
rect 366 61 379 62
rect 366 59 375 61
rect 377 59 379 61
rect 308 54 313 56
rect 277 45 290 46
rect 277 43 282 45
rect 284 43 290 45
rect 277 42 290 43
rect 222 31 224 32
rect 214 30 224 31
rect 226 30 227 32
rect 214 28 227 30
rect 214 26 216 28
rect 218 26 227 28
rect 214 25 227 26
rect 262 22 266 42
rect 284 37 298 38
rect 284 35 292 37
rect 294 35 298 37
rect 284 34 298 35
rect 308 52 309 54
rect 311 52 313 54
rect 308 47 313 52
rect 319 55 321 57
rect 323 55 324 57
rect 366 58 379 59
rect 319 54 324 55
rect 319 53 332 54
rect 319 51 329 53
rect 331 51 332 53
rect 319 50 332 51
rect 308 45 309 47
rect 311 45 313 47
rect 308 43 313 45
rect 284 25 289 34
rect 309 29 313 43
rect 309 27 310 29
rect 312 27 313 29
rect 309 23 313 27
rect 242 21 266 22
rect 242 19 244 21
rect 246 19 266 21
rect 242 18 266 19
rect 301 21 309 23
rect 311 21 313 23
rect 301 17 313 21
rect 333 37 339 39
rect 333 35 334 37
rect 336 35 339 37
rect 333 30 339 35
rect 326 29 339 30
rect 326 27 327 29
rect 329 27 339 29
rect 351 45 363 47
rect 351 43 352 45
rect 354 43 363 45
rect 351 42 363 43
rect 351 41 361 42
rect 359 40 361 41
rect 359 33 363 40
rect 375 37 379 58
rect 375 35 376 37
rect 378 35 379 37
rect 326 26 339 27
rect 375 25 379 35
rect 374 23 379 25
rect 374 21 375 23
rect 377 21 379 23
rect 374 19 379 21
rect 375 17 379 19
rect 386 61 399 62
rect 386 59 388 61
rect 390 59 399 61
rect 386 58 399 59
rect 386 25 390 58
rect 441 57 446 63
rect 441 55 442 57
rect 444 55 446 57
rect 441 54 446 55
rect 433 50 446 54
rect 453 61 466 62
rect 453 59 455 61
rect 457 59 466 61
rect 453 58 466 59
rect 402 42 414 47
rect 404 41 414 42
rect 404 40 406 41
rect 402 37 406 40
rect 402 35 403 37
rect 405 35 406 37
rect 402 33 406 35
rect 426 37 432 39
rect 426 35 429 37
rect 431 35 432 37
rect 426 30 432 35
rect 426 29 439 30
rect 426 27 434 29
rect 436 27 439 29
rect 426 26 439 27
rect 386 23 391 25
rect 386 21 388 23
rect 390 21 391 23
rect 386 19 391 21
rect 386 17 390 19
rect 453 29 457 58
rect 508 57 513 63
rect 508 55 509 57
rect 511 55 513 57
rect 508 54 513 55
rect 500 53 513 54
rect 500 51 501 53
rect 503 51 513 53
rect 500 50 513 51
rect 519 62 523 63
rect 519 58 532 62
rect 519 56 521 58
rect 519 51 523 56
rect 519 49 521 51
rect 469 44 481 47
rect 469 42 477 44
rect 479 42 481 44
rect 471 41 481 42
rect 471 40 473 41
rect 453 27 454 29
rect 456 27 457 29
rect 469 33 473 40
rect 453 25 457 27
rect 493 37 499 39
rect 493 35 496 37
rect 498 35 499 37
rect 493 30 499 35
rect 493 29 506 30
rect 493 27 502 29
rect 504 27 506 29
rect 493 26 506 27
rect 453 23 458 25
rect 453 21 455 23
rect 457 21 458 23
rect 453 19 458 21
rect 453 17 457 19
rect 519 45 523 49
rect 519 43 520 45
rect 522 43 523 45
rect 519 30 523 43
rect 551 46 555 55
rect 534 44 555 46
rect 534 42 548 44
rect 550 42 555 44
rect 561 54 577 55
rect 561 52 573 54
rect 575 52 577 54
rect 561 50 577 52
rect 519 28 524 30
rect 519 26 521 28
rect 523 26 524 28
rect 519 24 524 26
rect 534 37 555 38
rect 534 35 538 37
rect 540 35 555 37
rect 534 34 555 35
rect 551 25 555 34
rect 561 29 565 50
rect 609 57 621 63
rect 561 27 562 29
rect 564 27 565 29
rect 561 22 565 27
rect 600 32 605 39
rect 616 45 621 57
rect 616 43 617 45
rect 619 43 621 45
rect 616 41 621 43
rect 600 30 601 32
rect 603 31 605 32
rect 603 30 613 31
rect 600 25 613 30
rect 561 21 585 22
rect 561 19 581 21
rect 583 19 585 21
rect 561 18 585 19
rect -1 11 629 12
rect -1 9 6 11
rect 8 9 55 11
rect 57 9 65 11
rect 67 9 95 11
rect 97 9 148 11
rect 150 9 169 11
rect 171 9 179 11
rect 181 9 209 11
rect 211 9 262 11
rect 264 9 298 11
rect 300 9 308 11
rect 310 9 522 11
rect 524 9 563 11
rect 565 9 616 11
rect 618 9 629 11
rect -1 4 629 9
<< alu2 >>
rect 75 126 107 127
rect 75 124 76 126
rect 78 124 101 126
rect 103 124 107 126
rect 75 122 107 124
rect 147 126 221 127
rect 147 125 190 126
rect 147 123 148 125
rect 150 124 190 125
rect 192 124 215 126
rect 217 124 221 126
rect 150 123 221 124
rect 147 122 221 123
rect 308 125 329 126
rect 308 123 309 125
rect 311 123 326 125
rect 328 123 329 125
rect 308 122 329 123
rect 432 125 456 126
rect 432 123 433 125
rect 435 123 453 125
rect 455 123 456 125
rect 432 122 456 123
rect 500 125 564 126
rect 500 123 501 125
rect 503 123 561 125
rect 563 123 564 125
rect 500 122 564 123
rect 34 117 169 118
rect 34 115 35 117
rect 37 115 166 117
rect 168 115 169 117
rect 34 114 169 115
rect 374 117 405 118
rect 374 115 375 117
rect 377 115 402 117
rect 404 115 405 117
rect 374 114 405 115
rect 261 110 355 111
rect 261 108 262 110
rect 264 109 355 110
rect 264 108 351 109
rect 261 107 351 108
rect 353 107 355 109
rect 261 106 355 107
rect 475 110 522 111
rect 475 108 476 110
rect 478 109 522 110
rect 478 108 519 109
rect 475 107 519 108
rect 521 107 522 109
rect 475 106 522 107
rect 83 102 96 103
rect 83 100 84 102
rect 86 100 93 102
rect 95 100 96 102
rect 83 99 96 100
rect 197 102 210 103
rect 197 100 198 102
rect 200 100 207 102
rect 209 100 210 102
rect 197 99 210 100
rect 327 101 504 102
rect 327 99 328 101
rect 330 99 500 101
rect 502 99 504 101
rect 197 76 201 99
rect 327 98 504 99
rect 3 70 201 76
rect 3 55 8 70
rect 3 46 7 55
rect 328 53 505 54
rect 84 52 97 53
rect 84 50 85 52
rect 87 50 94 52
rect 96 50 97 52
rect 84 49 97 50
rect 198 52 211 53
rect 198 50 199 52
rect 201 50 208 52
rect 210 50 211 52
rect 328 51 329 53
rect 331 51 501 53
rect 503 51 505 53
rect 328 50 505 51
rect 198 49 211 50
rect 3 44 4 46
rect 6 44 7 46
rect 3 41 7 44
rect 262 45 356 46
rect 262 44 352 45
rect 262 42 263 44
rect 265 43 352 44
rect 354 43 356 45
rect 265 42 356 43
rect 262 41 356 42
rect 476 45 523 46
rect 476 44 520 45
rect 476 42 477 44
rect 479 43 520 44
rect 522 43 523 45
rect 479 42 523 43
rect 476 41 523 42
rect 35 37 170 38
rect 35 35 36 37
rect 38 35 167 37
rect 169 35 170 37
rect 35 34 170 35
rect 375 37 406 38
rect 375 35 376 37
rect 378 35 403 37
rect 405 35 406 37
rect 375 34 406 35
rect 76 28 108 30
rect 76 26 77 28
rect 79 26 102 28
rect 104 26 108 28
rect 76 25 108 26
rect 148 29 222 30
rect 148 27 149 29
rect 151 28 222 29
rect 151 27 191 28
rect 148 26 191 27
rect 193 26 216 28
rect 218 26 222 28
rect 309 29 330 30
rect 309 27 310 29
rect 312 27 327 29
rect 329 27 330 29
rect 309 26 330 27
rect 433 29 457 30
rect 433 27 434 29
rect 436 27 454 29
rect 456 27 457 29
rect 433 26 457 27
rect 501 29 565 30
rect 501 27 502 29
rect 504 27 562 29
rect 564 27 565 29
rect 501 26 565 27
rect 148 25 222 26
<< ptie >>
rect 3 143 9 145
rect 3 141 5 143
rect 7 141 9 143
rect 52 143 58 145
rect 52 141 54 143
rect 56 141 58 143
rect 3 139 9 141
rect 52 139 58 141
rect 92 143 98 145
rect 92 141 94 143
rect 96 141 98 143
rect 92 139 98 141
rect 166 143 172 145
rect 166 141 168 143
rect 170 141 172 143
rect 166 139 172 141
rect 206 143 212 145
rect 206 141 208 143
rect 210 141 212 143
rect 206 139 212 141
rect 305 143 311 145
rect 305 141 307 143
rect 309 141 311 143
rect 305 139 311 141
rect 519 143 525 145
rect 519 141 521 143
rect 523 141 525 143
rect 519 139 525 141
rect 613 143 619 145
rect 613 141 615 143
rect 617 141 619 143
rect 613 139 619 141
rect 4 11 10 13
rect 53 11 59 13
rect 4 9 6 11
rect 8 9 10 11
rect 4 7 10 9
rect 53 9 55 11
rect 57 9 59 11
rect 53 7 59 9
rect 93 11 99 13
rect 93 9 95 11
rect 97 9 99 11
rect 93 7 99 9
rect 167 11 173 13
rect 167 9 169 11
rect 171 9 173 11
rect 167 7 173 9
rect 207 11 213 13
rect 207 9 209 11
rect 211 9 213 11
rect 207 7 213 9
rect 306 11 312 13
rect 306 9 308 11
rect 310 9 312 11
rect 306 7 312 9
rect 520 11 526 13
rect 520 9 522 11
rect 524 9 526 11
rect 520 7 526 9
rect 614 11 620 13
rect 614 9 616 11
rect 618 9 620 11
rect 614 7 620 9
<< ntie >>
rect 3 83 9 85
rect 3 81 5 83
rect 7 81 9 83
rect 52 83 58 85
rect 3 79 9 81
rect 52 81 54 83
rect 56 81 58 83
rect 125 83 131 85
rect 52 79 58 81
rect 125 81 127 83
rect 129 81 131 83
rect 166 83 172 85
rect 125 79 131 81
rect 166 81 168 83
rect 170 81 172 83
rect 239 83 245 85
rect 166 79 172 81
rect 239 81 241 83
rect 243 81 245 83
rect 305 83 311 85
rect 239 79 245 81
rect 305 81 307 83
rect 309 81 311 83
rect 519 83 525 85
rect 305 79 311 81
rect 519 81 521 83
rect 523 81 525 83
rect 580 83 586 85
rect 519 79 525 81
rect 580 81 582 83
rect 584 81 586 83
rect 580 79 586 81
rect 4 71 10 73
rect 4 69 6 71
rect 8 69 10 71
rect 53 71 59 73
rect 4 67 10 69
rect 53 69 55 71
rect 57 69 59 71
rect 126 71 132 73
rect 53 67 59 69
rect 126 69 128 71
rect 130 69 132 71
rect 167 71 173 73
rect 126 67 132 69
rect 167 69 169 71
rect 171 69 173 71
rect 240 71 246 73
rect 167 67 173 69
rect 240 69 242 71
rect 244 69 246 71
rect 306 71 312 73
rect 240 67 246 69
rect 306 69 308 71
rect 310 69 312 71
rect 520 71 526 73
rect 306 67 312 69
rect 520 69 522 71
rect 524 69 526 71
rect 581 71 587 73
rect 520 67 526 69
rect 581 69 583 71
rect 585 69 587 71
rect 581 67 587 69
<< nmos >>
rect 9 122 11 131
rect 19 122 21 128
rect 29 122 31 128
rect 58 124 60 133
rect 71 124 73 135
rect 78 124 80 135
rect 98 122 100 131
rect 114 127 116 136
rect 124 127 126 136
rect 134 127 136 139
rect 141 127 143 139
rect 172 124 174 133
rect 185 124 187 135
rect 192 124 194 135
rect 212 122 214 131
rect 228 127 230 136
rect 238 127 240 136
rect 248 127 250 139
rect 255 127 257 139
rect 283 124 285 135
rect 290 124 292 135
rect 303 124 305 133
rect 325 128 327 134
rect 335 128 337 136
rect 342 128 344 136
rect 352 128 354 136
rect 359 128 361 136
rect 369 127 371 136
rect 392 127 394 136
rect 402 128 404 136
rect 409 128 411 136
rect 419 128 421 136
rect 426 128 428 136
rect 436 128 438 134
rect 459 127 461 136
rect 469 128 471 136
rect 476 128 478 136
rect 486 128 488 136
rect 493 128 495 136
rect 503 128 505 134
rect 525 122 527 131
rect 535 122 537 128
rect 545 122 547 128
rect 568 127 570 139
rect 575 127 577 139
rect 585 127 587 136
rect 595 127 597 136
rect 611 122 613 131
rect 10 21 12 30
rect 20 24 22 30
rect 30 24 32 30
rect 59 19 61 28
rect 72 17 74 28
rect 79 17 81 28
rect 99 21 101 30
rect 115 16 117 25
rect 125 16 127 25
rect 135 13 137 25
rect 142 13 144 25
rect 173 19 175 28
rect 186 17 188 28
rect 193 17 195 28
rect 213 21 215 30
rect 229 16 231 25
rect 239 16 241 25
rect 249 13 251 25
rect 256 13 258 25
rect 284 17 286 28
rect 291 17 293 28
rect 304 19 306 28
rect 326 18 328 24
rect 336 16 338 24
rect 343 16 345 24
rect 353 16 355 24
rect 360 16 362 24
rect 370 16 372 25
rect 393 16 395 25
rect 403 16 405 24
rect 410 16 412 24
rect 420 16 422 24
rect 427 16 429 24
rect 437 18 439 24
rect 460 16 462 25
rect 470 16 472 24
rect 477 16 479 24
rect 487 16 489 24
rect 494 16 496 24
rect 504 18 506 24
rect 526 21 528 30
rect 536 24 538 30
rect 546 24 548 30
rect 569 13 571 25
rect 576 13 578 25
rect 586 16 588 25
rect 596 16 598 25
rect 612 21 614 30
<< pmos >>
rect 9 92 11 110
rect 22 82 24 103
rect 29 82 31 103
rect 58 91 60 109
rect 68 89 70 102
rect 78 89 80 102
rect 106 82 108 109
rect 122 91 124 109
rect 132 91 134 109
rect 142 82 144 109
rect 172 91 174 109
rect 182 89 184 102
rect 192 89 194 102
rect 220 82 222 109
rect 236 91 238 109
rect 246 91 248 109
rect 256 82 258 109
rect 283 89 285 102
rect 293 89 295 102
rect 303 91 305 109
rect 325 102 327 110
rect 335 82 337 98
rect 342 82 344 98
rect 352 82 354 98
rect 359 82 361 98
rect 369 82 371 100
rect 392 82 394 100
rect 436 102 438 110
rect 402 82 404 98
rect 409 82 411 98
rect 419 82 421 98
rect 426 82 428 98
rect 459 82 461 100
rect 503 102 505 110
rect 469 82 471 98
rect 476 82 478 98
rect 486 82 488 98
rect 493 82 495 98
rect 525 92 527 110
rect 538 82 540 103
rect 545 82 547 103
rect 567 82 569 109
rect 577 91 579 109
rect 587 91 589 109
rect 603 82 605 109
rect 10 42 12 60
rect 23 49 25 70
rect 30 49 32 70
rect 59 43 61 61
rect 69 50 71 63
rect 79 50 81 63
rect 107 43 109 70
rect 123 43 125 61
rect 133 43 135 61
rect 143 43 145 70
rect 173 43 175 61
rect 183 50 185 63
rect 193 50 195 63
rect 221 43 223 70
rect 237 43 239 61
rect 247 43 249 61
rect 257 43 259 70
rect 284 50 286 63
rect 294 50 296 63
rect 304 43 306 61
rect 336 54 338 70
rect 343 54 345 70
rect 353 54 355 70
rect 360 54 362 70
rect 326 42 328 50
rect 370 52 372 70
rect 393 52 395 70
rect 403 54 405 70
rect 410 54 412 70
rect 420 54 422 70
rect 427 54 429 70
rect 460 52 462 70
rect 470 54 472 70
rect 477 54 479 70
rect 487 54 489 70
rect 494 54 496 70
rect 437 42 439 50
rect 504 42 506 50
rect 526 42 528 60
rect 539 49 541 70
rect 546 49 548 70
rect 568 43 570 70
rect 578 43 580 61
rect 588 43 590 61
rect 604 43 606 70
<< polyct0 >>
rect 11 115 13 117
rect 60 115 62 117
rect 130 115 132 117
rect 140 114 142 116
rect 174 115 176 117
rect 244 115 246 117
rect 254 114 256 116
rect 301 115 303 117
rect 350 121 352 123
rect 368 120 370 122
rect 393 120 395 122
rect 343 105 345 107
rect 411 121 413 123
rect 418 105 420 107
rect 460 120 462 122
rect 478 121 480 123
rect 485 105 487 107
rect 527 115 529 117
rect 569 114 571 116
rect 579 115 581 117
rect 12 35 14 37
rect 61 35 63 37
rect 131 35 133 37
rect 141 36 143 38
rect 175 35 177 37
rect 245 35 247 37
rect 255 36 257 38
rect 302 35 304 37
rect 344 45 346 47
rect 351 29 353 31
rect 419 45 421 47
rect 369 30 371 32
rect 394 30 396 32
rect 412 29 414 31
rect 486 45 488 47
rect 461 30 463 32
rect 479 29 481 31
rect 528 35 530 37
rect 570 36 572 38
rect 580 35 582 37
<< polyct1 >>
rect 21 115 23 117
rect 70 115 72 117
rect 31 108 33 110
rect 109 120 111 122
rect 80 107 82 109
rect 184 115 186 117
rect 93 107 95 109
rect 223 120 225 122
rect 194 107 196 109
rect 291 115 293 117
rect 207 107 209 109
rect 281 107 283 109
rect 333 115 335 117
rect 360 110 362 112
rect 401 110 403 112
rect 428 115 430 117
rect 320 95 322 97
rect 468 110 470 112
rect 495 115 497 117
rect 441 95 443 97
rect 537 115 539 117
rect 508 95 510 97
rect 600 120 602 122
rect 547 108 549 110
rect 616 107 618 109
rect 32 42 34 44
rect 22 35 24 37
rect 81 43 83 45
rect 94 43 96 45
rect 71 35 73 37
rect 195 43 197 45
rect 208 43 210 45
rect 282 43 284 45
rect 110 30 112 32
rect 185 35 187 37
rect 224 30 226 32
rect 321 55 323 57
rect 292 35 294 37
rect 442 55 444 57
rect 334 35 336 37
rect 361 40 363 42
rect 402 40 404 42
rect 509 55 511 57
rect 429 35 431 37
rect 469 40 471 42
rect 496 35 498 37
rect 548 42 550 44
rect 617 43 619 45
rect 538 35 540 37
rect 601 30 603 32
<< ndifct0 >>
rect 15 137 17 139
rect 34 137 36 139
rect 24 124 26 126
rect 83 131 85 133
rect 107 132 109 134
rect 93 124 95 126
rect 119 129 121 131
rect 197 131 199 133
rect 221 132 223 134
rect 207 124 209 126
rect 233 129 235 131
rect 278 131 280 133
rect 320 130 322 132
rect 330 130 332 132
rect 347 132 349 134
rect 364 132 366 134
rect 397 132 399 134
rect 414 132 416 134
rect 431 130 433 132
rect 441 130 443 132
rect 464 132 466 134
rect 481 132 483 134
rect 531 137 533 139
rect 498 130 500 132
rect 508 130 510 132
rect 550 137 552 139
rect 540 124 542 126
rect 590 129 592 131
rect 602 132 604 134
rect 616 124 618 126
rect 25 26 27 28
rect 16 13 18 15
rect 94 26 96 28
rect 84 19 86 21
rect 108 18 110 20
rect 35 13 37 15
rect 120 21 122 23
rect 208 26 210 28
rect 198 19 200 21
rect 222 18 224 20
rect 234 21 236 23
rect 279 19 281 21
rect 321 20 323 22
rect 331 20 333 22
rect 348 18 350 20
rect 365 18 367 20
rect 398 18 400 20
rect 415 18 417 20
rect 432 20 434 22
rect 442 20 444 22
rect 465 18 467 20
rect 482 18 484 20
rect 499 20 501 22
rect 509 20 511 22
rect 541 26 543 28
rect 532 13 534 15
rect 551 13 553 15
rect 591 21 593 23
rect 617 26 619 28
rect 603 18 605 20
<< ndifct1 >>
rect 64 141 66 143
rect 4 124 6 126
rect 147 141 149 143
rect 178 141 180 143
rect 53 129 55 131
rect 129 131 131 133
rect 261 141 263 143
rect 297 141 299 143
rect 167 129 169 131
rect 243 131 245 133
rect 308 129 310 131
rect 374 129 376 131
rect 387 129 389 131
rect 454 129 456 131
rect 562 141 564 143
rect 520 124 522 126
rect 580 131 582 133
rect 5 26 7 28
rect 54 21 56 23
rect 130 19 132 21
rect 65 9 67 11
rect 168 21 170 23
rect 148 9 150 11
rect 244 19 246 21
rect 179 9 181 11
rect 309 21 311 23
rect 262 9 264 11
rect 298 9 300 11
rect 375 21 377 23
rect 388 21 390 23
rect 455 21 457 23
rect 521 26 523 28
rect 581 19 583 21
rect 563 9 565 11
<< ntiect1 >>
rect 5 81 7 83
rect 54 81 56 83
rect 127 81 129 83
rect 168 81 170 83
rect 241 81 243 83
rect 307 81 309 83
rect 521 81 523 83
rect 582 81 584 83
rect 6 69 8 71
rect 55 69 57 71
rect 128 69 130 71
rect 169 69 171 71
rect 242 69 244 71
rect 308 69 310 71
rect 522 69 524 71
rect 583 69 585 71
<< ptiect1 >>
rect 5 141 7 143
rect 54 141 56 143
rect 94 141 96 143
rect 168 141 170 143
rect 208 141 210 143
rect 307 141 309 143
rect 521 141 523 143
rect 615 141 617 143
rect 6 9 8 11
rect 55 9 57 11
rect 95 9 97 11
rect 169 9 171 11
rect 209 9 211 11
rect 308 9 310 11
rect 522 9 524 11
rect 616 9 618 11
<< pdifct0 >>
rect 15 84 17 86
rect 34 91 36 93
rect 101 105 103 107
rect 63 93 65 95
rect 73 98 75 100
rect 73 91 75 93
rect 83 91 85 93
rect 111 91 113 93
rect 127 105 129 107
rect 127 98 129 100
rect 111 84 113 86
rect 147 90 149 92
rect 215 105 217 107
rect 177 93 179 95
rect 187 98 189 100
rect 187 91 189 93
rect 197 91 199 93
rect 225 91 227 93
rect 241 105 243 107
rect 241 98 243 100
rect 225 84 227 86
rect 261 90 263 92
rect 278 91 280 93
rect 288 98 290 100
rect 288 91 290 93
rect 298 93 300 95
rect 320 106 322 108
rect 330 84 332 86
rect 347 94 349 96
rect 364 84 366 86
rect 441 106 443 108
rect 397 84 399 86
rect 414 94 416 96
rect 431 84 433 86
rect 508 106 510 108
rect 464 84 466 86
rect 481 94 483 96
rect 498 84 500 86
rect 531 84 533 86
rect 550 91 552 93
rect 562 90 564 92
rect 582 105 584 107
rect 582 98 584 100
rect 598 91 600 93
rect 598 84 600 86
rect 608 105 610 107
rect 16 66 18 68
rect 35 59 37 61
rect 64 57 66 59
rect 74 59 76 61
rect 74 52 76 54
rect 84 59 86 61
rect 102 45 104 47
rect 112 66 114 68
rect 112 59 114 61
rect 128 52 130 54
rect 128 45 130 47
rect 148 60 150 62
rect 178 57 180 59
rect 188 59 190 61
rect 188 52 190 54
rect 198 59 200 61
rect 216 45 218 47
rect 226 66 228 68
rect 226 59 228 61
rect 242 52 244 54
rect 242 45 244 47
rect 331 66 333 68
rect 262 60 264 62
rect 279 59 281 61
rect 289 59 291 61
rect 289 52 291 54
rect 299 57 301 59
rect 348 56 350 58
rect 365 66 367 68
rect 321 44 323 46
rect 398 66 400 68
rect 415 56 417 58
rect 432 66 434 68
rect 465 66 467 68
rect 482 56 484 58
rect 499 66 501 68
rect 532 66 534 68
rect 442 44 444 46
rect 509 44 511 46
rect 551 59 553 61
rect 563 60 565 62
rect 599 66 601 68
rect 583 52 585 54
rect 583 45 585 47
rect 599 59 601 61
rect 609 45 611 47
<< pdifct1 >>
rect 4 101 6 103
rect 4 94 6 96
rect 53 105 55 107
rect 53 98 55 100
rect 137 98 139 100
rect 167 105 169 107
rect 167 98 169 100
rect 251 98 253 100
rect 308 105 310 107
rect 308 98 310 100
rect 374 91 376 93
rect 387 91 389 93
rect 454 91 456 93
rect 520 101 522 103
rect 520 94 522 96
rect 572 98 574 100
rect 5 56 7 58
rect 5 49 7 51
rect 54 52 56 54
rect 54 45 56 47
rect 138 52 140 54
rect 168 52 170 54
rect 168 45 170 47
rect 252 52 254 54
rect 309 52 311 54
rect 309 45 311 47
rect 375 59 377 61
rect 388 59 390 61
rect 455 59 457 61
rect 521 56 523 58
rect 521 49 523 51
rect 573 52 575 54
<< alu0 >>
rect 13 139 19 140
rect 13 137 15 139
rect 17 137 19 139
rect 13 136 19 137
rect 32 139 38 140
rect 32 137 34 139
rect 36 137 38 139
rect 32 136 38 137
rect 105 134 111 140
rect 67 133 87 134
rect 67 131 83 133
rect 85 131 87 133
rect 105 132 107 134
rect 109 132 111 134
rect 105 131 111 132
rect 118 131 122 133
rect 67 130 87 131
rect 10 126 28 127
rect 10 124 24 126
rect 26 124 28 126
rect 10 123 28 124
rect 10 117 14 123
rect 10 115 11 117
rect 13 115 14 117
rect 6 94 7 105
rect 10 102 14 115
rect 29 110 35 111
rect 55 127 56 129
rect 67 126 71 130
rect 118 129 119 131
rect 121 129 122 131
rect 59 122 71 126
rect 59 117 63 122
rect 59 115 60 117
rect 62 115 63 117
rect 10 98 25 102
rect 21 94 25 98
rect 59 103 63 115
rect 92 126 96 128
rect 92 124 93 126
rect 95 124 96 126
rect 92 118 96 124
rect 118 126 122 129
rect 118 122 142 126
rect 92 114 103 118
rect 59 100 76 103
rect 59 99 73 100
rect 72 98 73 99
rect 75 98 76 100
rect 61 95 67 96
rect 21 93 38 94
rect 21 91 34 93
rect 36 91 38 93
rect 21 90 38 91
rect 61 93 63 95
rect 65 93 67 95
rect 13 86 19 87
rect 13 84 15 86
rect 17 84 19 86
rect 61 84 67 93
rect 72 93 76 98
rect 99 108 103 114
rect 138 118 142 122
rect 118 117 134 118
rect 118 115 130 117
rect 132 115 134 117
rect 118 114 134 115
rect 138 116 143 118
rect 138 114 140 116
rect 142 114 143 116
rect 118 108 122 114
rect 138 112 143 114
rect 138 110 142 112
rect 99 107 122 108
rect 99 105 101 107
rect 103 105 122 107
rect 99 104 122 105
rect 72 91 73 93
rect 75 91 76 93
rect 72 89 76 91
rect 81 93 87 94
rect 81 91 83 93
rect 85 91 87 93
rect 81 84 87 91
rect 110 93 114 95
rect 110 91 111 93
rect 113 91 114 93
rect 110 86 114 91
rect 118 93 122 104
rect 126 107 142 110
rect 126 105 127 107
rect 129 106 142 107
rect 129 105 130 106
rect 126 100 130 105
rect 126 98 127 100
rect 129 98 130 100
rect 126 96 130 98
rect 219 134 225 140
rect 181 133 201 134
rect 181 131 197 133
rect 199 131 201 133
rect 219 132 221 134
rect 223 132 225 134
rect 219 131 225 132
rect 232 131 236 133
rect 181 130 201 131
rect 169 127 170 129
rect 181 126 185 130
rect 232 129 233 131
rect 235 129 236 131
rect 276 133 296 134
rect 276 131 278 133
rect 280 131 296 133
rect 276 130 296 131
rect 173 122 185 126
rect 173 117 177 122
rect 173 115 174 117
rect 176 115 177 117
rect 173 103 177 115
rect 206 126 210 128
rect 206 124 207 126
rect 209 124 210 126
rect 206 118 210 124
rect 232 126 236 129
rect 232 122 256 126
rect 206 114 217 118
rect 173 100 190 103
rect 173 99 187 100
rect 186 98 187 99
rect 189 98 190 100
rect 175 95 181 96
rect 175 93 177 95
rect 179 93 181 95
rect 118 92 151 93
rect 118 90 147 92
rect 149 90 151 92
rect 118 89 151 90
rect 110 84 111 86
rect 113 84 114 86
rect 175 84 181 93
rect 186 93 190 98
rect 213 108 217 114
rect 252 118 256 122
rect 232 117 248 118
rect 232 115 244 117
rect 246 115 248 117
rect 232 114 248 115
rect 252 116 257 118
rect 252 114 254 116
rect 256 114 257 116
rect 232 108 236 114
rect 252 112 257 114
rect 252 110 256 112
rect 213 107 236 108
rect 213 105 215 107
rect 217 105 236 107
rect 213 104 236 105
rect 186 91 187 93
rect 189 91 190 93
rect 186 89 190 91
rect 195 93 201 94
rect 195 91 197 93
rect 199 91 201 93
rect 195 84 201 91
rect 224 93 228 95
rect 224 91 225 93
rect 227 91 228 93
rect 224 86 228 91
rect 232 93 236 104
rect 240 107 256 110
rect 240 105 241 107
rect 243 106 256 107
rect 292 126 296 130
rect 307 127 308 129
rect 292 122 304 126
rect 300 117 304 122
rect 300 115 301 117
rect 303 115 304 117
rect 243 105 244 106
rect 240 100 244 105
rect 240 98 241 100
rect 243 98 244 100
rect 240 96 244 98
rect 300 103 304 115
rect 287 100 304 103
rect 287 98 288 100
rect 290 99 304 100
rect 318 132 324 133
rect 318 130 320 132
rect 322 130 324 132
rect 318 129 324 130
rect 328 132 334 140
rect 328 130 330 132
rect 332 130 334 132
rect 345 134 360 135
rect 345 132 347 134
rect 349 132 360 134
rect 345 131 360 132
rect 328 129 334 130
rect 318 109 322 129
rect 356 126 360 131
rect 363 134 367 140
rect 363 132 364 134
rect 366 132 367 134
rect 363 130 367 132
rect 342 123 353 125
rect 342 121 350 123
rect 352 121 353 123
rect 356 124 370 126
rect 356 122 371 124
rect 342 119 353 121
rect 366 120 368 122
rect 370 120 371 122
rect 342 109 346 119
rect 366 118 371 120
rect 318 108 346 109
rect 318 106 320 108
rect 322 107 346 108
rect 322 106 343 107
rect 318 105 343 106
rect 345 105 346 107
rect 362 108 363 114
rect 342 103 346 105
rect 290 98 291 99
rect 276 93 282 94
rect 232 92 265 93
rect 232 90 261 92
rect 263 90 265 92
rect 232 89 265 90
rect 276 91 278 93
rect 280 91 282 93
rect 224 84 225 86
rect 227 84 228 86
rect 276 84 282 91
rect 287 93 291 98
rect 366 101 370 118
rect 354 97 370 101
rect 287 91 288 93
rect 290 91 291 93
rect 287 89 291 91
rect 296 95 302 96
rect 296 93 298 95
rect 300 93 302 95
rect 296 84 302 93
rect 345 96 358 97
rect 345 94 347 96
rect 349 94 358 96
rect 345 93 358 94
rect 396 134 400 140
rect 396 132 397 134
rect 399 132 400 134
rect 396 130 400 132
rect 403 134 418 135
rect 403 132 414 134
rect 416 132 418 134
rect 403 131 418 132
rect 429 132 435 140
rect 463 134 467 140
rect 403 126 407 131
rect 429 130 431 132
rect 433 130 435 132
rect 429 129 435 130
rect 439 132 445 133
rect 439 130 441 132
rect 443 130 445 132
rect 439 129 445 130
rect 393 124 407 126
rect 392 122 407 124
rect 410 123 421 125
rect 392 120 393 122
rect 395 120 397 122
rect 392 118 397 120
rect 410 121 411 123
rect 413 121 421 123
rect 410 119 421 121
rect 393 101 397 118
rect 400 108 401 114
rect 417 109 421 119
rect 441 109 445 129
rect 417 108 445 109
rect 417 107 441 108
rect 417 105 418 107
rect 420 106 441 107
rect 443 106 445 108
rect 420 105 445 106
rect 463 132 464 134
rect 466 132 467 134
rect 463 130 467 132
rect 470 134 485 135
rect 470 132 481 134
rect 483 132 485 134
rect 470 131 485 132
rect 496 132 502 140
rect 529 139 535 140
rect 529 137 531 139
rect 533 137 535 139
rect 529 136 535 137
rect 548 139 554 140
rect 548 137 550 139
rect 552 137 554 139
rect 548 136 554 137
rect 600 134 606 140
rect 470 126 474 131
rect 496 130 498 132
rect 500 130 502 132
rect 496 129 502 130
rect 506 132 512 133
rect 506 130 508 132
rect 510 130 512 132
rect 506 129 512 130
rect 460 124 474 126
rect 417 103 421 105
rect 393 97 409 101
rect 405 96 418 97
rect 405 94 414 96
rect 416 94 418 96
rect 405 93 418 94
rect 459 122 474 124
rect 477 123 488 125
rect 459 120 460 122
rect 462 120 464 122
rect 459 118 464 120
rect 477 121 478 123
rect 480 121 488 123
rect 477 119 488 121
rect 460 101 464 118
rect 467 108 468 114
rect 484 109 488 119
rect 508 109 512 129
rect 589 131 593 133
rect 600 132 602 134
rect 604 132 606 134
rect 600 131 606 132
rect 484 108 512 109
rect 484 107 508 108
rect 484 105 485 107
rect 487 106 508 107
rect 510 106 512 108
rect 487 105 512 106
rect 526 126 544 127
rect 526 124 540 126
rect 542 124 544 126
rect 526 123 544 124
rect 484 103 488 105
rect 526 117 530 123
rect 526 115 527 117
rect 529 115 530 117
rect 460 97 476 101
rect 472 96 485 97
rect 472 94 481 96
rect 483 94 485 96
rect 472 93 485 94
rect 522 94 523 105
rect 526 102 530 115
rect 589 129 590 131
rect 592 129 593 131
rect 589 126 593 129
rect 545 110 551 111
rect 526 98 541 102
rect 537 94 541 98
rect 569 122 593 126
rect 569 118 573 122
rect 615 126 619 128
rect 615 124 616 126
rect 618 124 619 126
rect 568 116 573 118
rect 568 114 569 116
rect 571 114 573 116
rect 577 117 593 118
rect 577 115 579 117
rect 581 115 593 117
rect 577 114 593 115
rect 568 112 573 114
rect 569 110 573 112
rect 569 107 585 110
rect 569 106 582 107
rect 581 105 582 106
rect 584 105 585 107
rect 581 100 585 105
rect 581 98 582 100
rect 584 98 585 100
rect 581 96 585 98
rect 589 108 593 114
rect 615 118 619 124
rect 608 114 619 118
rect 608 108 612 114
rect 589 107 612 108
rect 589 105 608 107
rect 610 105 612 107
rect 589 104 612 105
rect 537 93 554 94
rect 589 93 593 104
rect 537 91 550 93
rect 552 91 554 93
rect 537 90 554 91
rect 560 92 593 93
rect 560 90 562 92
rect 564 90 593 92
rect 560 89 593 90
rect 597 93 601 95
rect 597 91 598 93
rect 600 91 601 93
rect 329 86 333 88
rect 329 84 330 86
rect 332 84 333 86
rect 362 86 368 87
rect 362 84 364 86
rect 366 84 368 86
rect 395 86 401 87
rect 395 84 397 86
rect 399 84 401 86
rect 430 86 434 88
rect 430 84 431 86
rect 433 84 434 86
rect 462 86 468 87
rect 462 84 464 86
rect 466 84 468 86
rect 497 86 501 88
rect 497 84 498 86
rect 500 84 501 86
rect 529 86 535 87
rect 529 84 531 86
rect 533 84 535 86
rect 597 86 601 91
rect 597 84 598 86
rect 600 84 601 86
rect 14 66 16 68
rect 18 66 20 68
rect 14 65 20 66
rect 22 61 39 62
rect 22 59 35 61
rect 37 59 39 61
rect 22 58 39 59
rect 62 59 68 68
rect 7 47 8 58
rect 22 54 26 58
rect 62 57 64 59
rect 66 57 68 59
rect 62 56 68 57
rect 73 61 77 63
rect 73 59 74 61
rect 76 59 77 61
rect 11 50 26 54
rect 73 54 77 59
rect 82 61 88 68
rect 111 66 112 68
rect 114 66 115 68
rect 82 59 84 61
rect 86 59 88 61
rect 82 58 88 59
rect 111 61 115 66
rect 111 59 112 61
rect 114 59 115 61
rect 111 57 115 59
rect 119 62 152 63
rect 119 60 148 62
rect 150 60 152 62
rect 119 59 152 60
rect 176 59 182 68
rect 73 53 74 54
rect 11 37 15 50
rect 60 52 74 53
rect 76 52 77 54
rect 60 49 77 52
rect 30 41 36 42
rect 11 35 12 37
rect 14 35 15 37
rect 11 29 15 35
rect 11 28 29 29
rect 11 26 25 28
rect 27 26 29 28
rect 11 25 29 26
rect 60 37 64 49
rect 119 48 123 59
rect 176 57 178 59
rect 180 57 182 59
rect 176 56 182 57
rect 187 61 191 63
rect 187 59 188 61
rect 190 59 191 61
rect 100 47 123 48
rect 100 45 102 47
rect 104 45 123 47
rect 100 44 123 45
rect 100 38 104 44
rect 60 35 61 37
rect 63 35 64 37
rect 60 30 64 35
rect 60 26 72 30
rect 56 23 57 25
rect 68 22 72 26
rect 93 34 104 38
rect 93 28 97 34
rect 119 38 123 44
rect 127 54 131 56
rect 127 52 128 54
rect 130 52 131 54
rect 127 47 131 52
rect 127 45 128 47
rect 130 46 131 47
rect 130 45 143 46
rect 127 42 143 45
rect 139 40 143 42
rect 139 38 144 40
rect 119 37 135 38
rect 119 35 131 37
rect 133 35 135 37
rect 119 34 135 35
rect 139 36 141 38
rect 143 36 144 38
rect 139 34 144 36
rect 93 26 94 28
rect 96 26 97 28
rect 93 24 97 26
rect 139 30 143 34
rect 119 26 143 30
rect 119 23 123 26
rect 68 21 88 22
rect 119 21 120 23
rect 122 21 123 23
rect 68 19 84 21
rect 86 19 88 21
rect 68 18 88 19
rect 106 20 112 21
rect 106 18 108 20
rect 110 18 112 20
rect 119 19 123 21
rect 187 54 191 59
rect 196 61 202 68
rect 225 66 226 68
rect 228 66 229 68
rect 196 59 198 61
rect 200 59 202 61
rect 196 58 202 59
rect 225 61 229 66
rect 225 59 226 61
rect 228 59 229 61
rect 225 57 229 59
rect 233 62 266 63
rect 233 60 262 62
rect 264 60 266 62
rect 233 59 266 60
rect 277 61 283 68
rect 277 59 279 61
rect 281 59 283 61
rect 187 53 188 54
rect 174 52 188 53
rect 190 52 191 54
rect 174 49 191 52
rect 174 37 178 49
rect 233 48 237 59
rect 277 58 283 59
rect 288 61 292 63
rect 288 59 289 61
rect 291 59 292 61
rect 214 47 237 48
rect 214 45 216 47
rect 218 45 237 47
rect 214 44 237 45
rect 214 38 218 44
rect 174 35 175 37
rect 177 35 178 37
rect 174 30 178 35
rect 174 26 186 30
rect 170 23 171 25
rect 14 15 20 16
rect 14 13 16 15
rect 18 13 20 15
rect 14 12 20 13
rect 33 15 39 16
rect 33 13 35 15
rect 37 13 39 15
rect 33 12 39 13
rect 106 12 112 18
rect 182 22 186 26
rect 207 34 218 38
rect 207 28 211 34
rect 233 38 237 44
rect 241 54 245 56
rect 241 52 242 54
rect 244 52 245 54
rect 241 47 245 52
rect 241 45 242 47
rect 244 46 245 47
rect 244 45 257 46
rect 241 42 257 45
rect 253 40 257 42
rect 288 54 292 59
rect 297 59 303 68
rect 330 66 331 68
rect 333 66 334 68
rect 330 64 334 66
rect 363 66 365 68
rect 367 66 369 68
rect 363 65 369 66
rect 396 66 398 68
rect 400 66 402 68
rect 396 65 402 66
rect 431 66 432 68
rect 434 66 435 68
rect 431 64 435 66
rect 463 66 465 68
rect 467 66 469 68
rect 463 65 469 66
rect 498 66 499 68
rect 501 66 502 68
rect 498 64 502 66
rect 530 66 532 68
rect 534 66 536 68
rect 530 65 536 66
rect 598 66 599 68
rect 601 66 602 68
rect 297 57 299 59
rect 301 57 303 59
rect 297 56 303 57
rect 288 52 289 54
rect 291 53 292 54
rect 291 52 305 53
rect 288 49 305 52
rect 253 38 258 40
rect 233 37 249 38
rect 233 35 245 37
rect 247 35 249 37
rect 233 34 249 35
rect 253 36 255 38
rect 257 36 258 38
rect 253 34 258 36
rect 207 26 208 28
rect 210 26 211 28
rect 207 24 211 26
rect 253 30 257 34
rect 233 26 257 30
rect 233 23 237 26
rect 182 21 202 22
rect 233 21 234 23
rect 236 21 237 23
rect 301 37 305 49
rect 346 58 359 59
rect 346 56 348 58
rect 350 56 359 58
rect 346 55 359 56
rect 355 51 371 55
rect 343 47 347 49
rect 301 35 302 37
rect 304 35 305 37
rect 301 30 305 35
rect 293 26 305 30
rect 293 22 297 26
rect 308 23 309 25
rect 182 19 198 21
rect 200 19 202 21
rect 182 18 202 19
rect 220 20 226 21
rect 220 18 222 20
rect 224 18 226 20
rect 233 19 237 21
rect 277 21 297 22
rect 277 19 279 21
rect 281 19 297 21
rect 277 18 297 19
rect 220 12 226 18
rect 319 46 344 47
rect 319 44 321 46
rect 323 45 344 46
rect 346 45 347 47
rect 323 44 347 45
rect 319 43 347 44
rect 319 23 323 43
rect 343 33 347 43
rect 363 38 364 44
rect 367 34 371 51
rect 343 31 354 33
rect 343 29 351 31
rect 353 29 354 31
rect 367 32 372 34
rect 367 30 369 32
rect 371 30 372 32
rect 343 27 354 29
rect 357 28 372 30
rect 357 26 371 28
rect 319 22 325 23
rect 319 20 321 22
rect 323 20 325 22
rect 319 19 325 20
rect 329 22 335 23
rect 329 20 331 22
rect 333 20 335 22
rect 357 21 361 26
rect 329 12 335 20
rect 346 20 361 21
rect 346 18 348 20
rect 350 18 361 20
rect 346 17 361 18
rect 364 20 368 22
rect 364 18 365 20
rect 367 18 368 20
rect 364 12 368 18
rect 406 58 419 59
rect 406 56 415 58
rect 417 56 419 58
rect 406 55 419 56
rect 394 51 410 55
rect 394 34 398 51
rect 473 58 486 59
rect 418 47 422 49
rect 401 38 402 44
rect 418 45 419 47
rect 421 46 446 47
rect 421 45 442 46
rect 418 44 442 45
rect 444 44 446 46
rect 418 43 446 44
rect 393 32 398 34
rect 418 33 422 43
rect 393 30 394 32
rect 396 30 398 32
rect 411 31 422 33
rect 393 28 408 30
rect 394 26 408 28
rect 411 29 412 31
rect 414 29 422 31
rect 411 27 422 29
rect 397 20 401 22
rect 397 18 398 20
rect 400 18 401 20
rect 397 12 401 18
rect 404 21 408 26
rect 442 23 446 43
rect 430 22 436 23
rect 404 20 419 21
rect 404 18 415 20
rect 417 18 419 20
rect 404 17 419 18
rect 430 20 432 22
rect 434 20 436 22
rect 430 12 436 20
rect 440 22 446 23
rect 440 20 442 22
rect 444 20 446 22
rect 440 19 446 20
rect 473 56 482 58
rect 484 56 486 58
rect 473 55 486 56
rect 461 51 477 55
rect 461 34 465 51
rect 561 62 594 63
rect 538 61 555 62
rect 538 59 551 61
rect 553 59 555 61
rect 561 60 563 62
rect 565 60 594 62
rect 561 59 594 60
rect 538 58 555 59
rect 485 47 489 49
rect 468 38 469 44
rect 485 45 486 47
rect 488 46 513 47
rect 488 45 509 46
rect 485 44 509 45
rect 511 44 513 46
rect 485 43 513 44
rect 460 32 465 34
rect 485 33 489 43
rect 460 30 461 32
rect 463 30 465 32
rect 478 31 489 33
rect 460 28 475 30
rect 461 26 475 28
rect 478 29 479 31
rect 481 29 489 31
rect 478 27 489 29
rect 464 20 468 22
rect 464 18 465 20
rect 467 18 468 20
rect 464 12 468 18
rect 471 21 475 26
rect 509 23 513 43
rect 523 47 524 58
rect 538 54 542 58
rect 527 50 542 54
rect 527 37 531 50
rect 582 54 586 56
rect 582 52 583 54
rect 585 52 586 54
rect 546 41 552 42
rect 527 35 528 37
rect 530 35 531 37
rect 527 29 531 35
rect 527 28 545 29
rect 527 26 541 28
rect 543 26 545 28
rect 527 25 545 26
rect 582 47 586 52
rect 582 46 583 47
rect 570 45 583 46
rect 585 45 586 47
rect 570 42 586 45
rect 590 48 594 59
rect 598 61 602 66
rect 598 59 599 61
rect 601 59 602 61
rect 598 57 602 59
rect 590 47 613 48
rect 590 45 609 47
rect 611 45 613 47
rect 590 44 613 45
rect 570 40 574 42
rect 569 38 574 40
rect 590 38 594 44
rect 569 36 570 38
rect 572 36 574 38
rect 569 34 574 36
rect 578 37 594 38
rect 578 35 580 37
rect 582 35 594 37
rect 578 34 594 35
rect 497 22 503 23
rect 471 20 486 21
rect 471 18 482 20
rect 484 18 486 20
rect 471 17 486 18
rect 497 20 499 22
rect 501 20 503 22
rect 497 12 503 20
rect 507 22 513 23
rect 507 20 509 22
rect 511 20 513 22
rect 507 19 513 20
rect 570 30 574 34
rect 609 38 613 44
rect 609 34 620 38
rect 570 26 594 30
rect 590 23 594 26
rect 616 28 620 34
rect 616 26 617 28
rect 619 26 620 28
rect 616 24 620 26
rect 590 21 591 23
rect 593 21 594 23
rect 590 19 594 21
rect 601 20 607 21
rect 601 18 603 20
rect 605 18 607 20
rect 530 15 536 16
rect 530 13 532 15
rect 534 13 536 15
rect 530 12 536 13
rect 549 15 555 16
rect 549 13 551 15
rect 553 13 555 15
rect 549 12 555 13
rect 601 12 607 18
<< via1 >>
rect 35 115 37 117
rect 76 124 78 126
rect 101 124 103 126
rect 84 100 86 102
rect 148 123 150 125
rect 93 100 95 102
rect 166 115 168 117
rect 190 124 192 126
rect 215 124 217 126
rect 198 100 200 102
rect 207 100 209 102
rect 262 108 264 110
rect 309 123 311 125
rect 326 123 328 125
rect 351 107 353 109
rect 328 99 330 101
rect 375 115 377 117
rect 402 115 404 117
rect 433 123 435 125
rect 453 123 455 125
rect 476 108 478 110
rect 501 123 503 125
rect 519 107 521 109
rect 500 99 502 101
rect 561 123 563 125
rect 4 44 6 46
rect 85 50 87 52
rect 36 35 38 37
rect 94 50 96 52
rect 77 26 79 28
rect 102 26 104 28
rect 149 27 151 29
rect 199 50 201 52
rect 167 35 169 37
rect 208 50 210 52
rect 191 26 193 28
rect 263 42 265 44
rect 216 26 218 28
rect 329 51 331 53
rect 310 27 312 29
rect 327 27 329 29
rect 352 43 354 45
rect 376 35 378 37
rect 403 35 405 37
rect 434 27 436 29
rect 501 51 503 53
rect 477 42 479 44
rect 454 27 456 29
rect 502 27 504 29
rect 520 43 522 45
rect 562 27 564 29
<< labels >>
rlabel alu1 122 8 122 8 6 vss
rlabel alu1 122 72 122 72 6 vdd
rlabel alu1 70 72 70 72 6 vdd
rlabel alu1 70 8 70 8 6 vss
rlabel alu1 236 8 236 8 6 vss
rlabel alu1 236 72 236 72 6 vdd
rlabel alu1 264 32 264 32 1 sum
rlabel alu1 184 72 184 72 6 vdd
rlabel alu1 184 8 184 8 6 vss
rlabel alu1 21 8 21 8 6 vss
rlabel alu1 21 72 21 72 6 vdd
rlabel alu1 70 35 70 35 1 a
rlabel via1 85 50 85 50 1 b
rlabel via1 201 51 201 51 1 cin
rlabel alu1 5 38 5 38 1 cout
rlabel alu1 295 8 295 8 4 vss
rlabel alu1 295 36 295 36 4 a
rlabel alu1 287 32 287 32 4 a
rlabel alu1 287 44 287 44 4 b
rlabel alu1 295 72 295 72 4 vdd
rlabel alu1 279 52 279 52 4 b
rlabel alu1 388 36 388 36 6 z
rlabel alu1 396 60 396 60 6 z
rlabel alu1 416 8 416 8 6 vss
rlabel alu1 416 72 416 72 6 vdd
rlabel via1 353 44 353 44 4 a0
rlabel alu1 361 40 361 40 4 a0
rlabel alu1 349 8 349 8 4 vss
rlabel alu1 337 36 337 36 4 a1
rlabel alu1 349 72 349 72 4 vdd
rlabel alu1 329 28 329 28 4 a1
rlabel alu1 483 8 483 8 6 vss
rlabel alu1 483 72 483 72 6 vdd
rlabel alu1 475 43 475 43 1 a2
rlabel alu1 471 38 471 38 1 a2
rlabel alu1 494 36 494 36 1 a3
rlabel alu1 499 27 499 27 1 a3
rlabel via1 503 52 503 52 1 s1
rlabel alu1 511 60 511 60 1 s1
rlabel via1 329 52 329 52 1 s1
rlabel alu1 321 60 321 60 1 s1
rlabel alu1 444 60 444 60 1 s0
rlabel alu1 537 8 537 8 6 vss
rlabel alu1 537 72 537 72 6 vdd
rlabel alu1 553 52 553 52 6 b
rlabel alu1 553 28 553 28 6 a
rlabel alu1 537 44 537 44 6 b
rlabel alu1 545 44 545 44 6 b
rlabel alu1 545 36 545 36 6 a
rlabel alu1 537 36 537 36 6 a
rlabel alu1 611 28 611 28 4 a
rlabel alu1 619 52 619 52 4 b
rlabel alu1 611 60 611 60 4 b
rlabel alu1 603 32 603 32 4 a
rlabel alu1 591 8 591 8 4 vss
rlabel alu1 591 72 591 72 4 vdd
rlabel alu1 121 144 121 144 8 vss
rlabel alu1 121 80 121 80 8 vdd
rlabel alu1 69 80 69 80 8 vdd
rlabel alu1 69 144 69 144 8 vss
rlabel alu1 235 144 235 144 8 vss
rlabel alu1 235 80 235 80 8 vdd
rlabel alu1 263 120 263 120 5 sum
rlabel alu1 183 80 183 80 8 vdd
rlabel alu1 183 144 183 144 8 vss
rlabel alu1 20 144 20 144 8 vss
rlabel alu1 20 80 20 80 8 vdd
rlabel alu1 69 117 69 117 5 a
rlabel via1 84 102 84 102 5 b
rlabel via1 200 101 200 101 5 cin
rlabel alu1 4 114 4 114 5 cout
rlabel alu1 294 144 294 144 2 vss
rlabel alu1 294 116 294 116 2 a
rlabel alu1 286 120 286 120 2 a
rlabel alu1 286 108 286 108 2 b
rlabel alu1 294 80 294 80 2 vdd
rlabel alu1 278 100 278 100 2 b
rlabel alu1 387 116 387 116 8 z
rlabel alu1 395 92 395 92 8 z
rlabel alu1 415 144 415 144 8 vss
rlabel alu1 415 80 415 80 8 vdd
rlabel via1 352 108 352 108 2 a0
rlabel alu1 360 112 360 112 2 a0
rlabel alu1 348 144 348 144 2 vss
rlabel alu1 336 116 336 116 2 a1
rlabel alu1 348 80 348 80 2 vdd
rlabel alu1 328 124 328 124 2 a1
rlabel alu1 482 144 482 144 8 vss
rlabel alu1 482 80 482 80 8 vdd
rlabel alu1 474 109 474 109 5 a2
rlabel alu1 470 114 470 114 5 a2
rlabel alu1 493 116 493 116 5 a3
rlabel alu1 498 125 498 125 5 a3
rlabel via1 502 100 502 100 5 s1
rlabel alu1 510 92 510 92 5 s1
rlabel via1 328 100 328 100 5 s1
rlabel alu1 320 92 320 92 5 s1
rlabel alu1 443 92 443 92 5 s0
rlabel alu1 536 144 536 144 8 vss
rlabel alu1 536 80 536 80 8 vdd
rlabel alu1 552 100 552 100 8 b
rlabel alu1 552 124 552 124 8 a
rlabel alu1 536 108 536 108 8 b
rlabel alu1 544 108 544 108 8 b
rlabel alu1 544 116 544 116 8 a
rlabel alu1 536 116 536 116 8 a
rlabel alu1 610 124 610 124 2 a
rlabel alu1 618 100 618 100 2 b
rlabel alu1 610 92 610 92 2 b
rlabel alu1 602 120 602 120 2 a
rlabel alu1 590 144 590 144 2 vss
rlabel alu1 590 80 590 80 2 vdd
<< end >>
