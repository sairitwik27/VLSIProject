magic
tech scmos
timestamp 1608824715
<< ab >>
rect 5 5 85 293
rect 87 5 190 293
rect 192 5 255 293
<< nwell >>
rect 0 181 260 261
rect 0 37 260 117
<< pwell >>
rect 0 261 260 298
rect 0 117 260 181
rect 0 0 260 37
<< poly >>
rect 14 276 16 281
rect 24 273 26 278
rect 34 273 36 278
rect 54 278 56 282
rect 67 280 69 285
rect 74 280 76 285
rect 98 289 123 291
rect 98 281 100 289
rect 111 281 113 285
rect 121 281 123 289
rect 131 284 133 289
rect 138 284 140 289
rect 95 279 100 281
rect 95 276 97 279
rect 14 264 16 267
rect 24 264 26 267
rect 14 262 20 264
rect 14 260 16 262
rect 18 260 20 262
rect 14 258 20 260
rect 24 262 30 264
rect 24 260 26 262
rect 28 260 30 262
rect 24 258 30 260
rect 14 255 16 258
rect 27 248 29 258
rect 34 257 36 267
rect 54 264 56 269
rect 67 264 69 269
rect 54 262 60 264
rect 54 260 56 262
rect 58 260 60 262
rect 54 258 60 260
rect 64 262 70 264
rect 64 260 66 262
rect 68 260 70 262
rect 64 258 70 260
rect 34 255 40 257
rect 34 253 36 255
rect 38 253 40 255
rect 54 254 56 258
rect 34 251 40 253
rect 34 248 36 251
rect 14 232 16 237
rect 64 247 66 258
rect 74 256 76 269
rect 159 278 161 282
rect 172 280 174 285
rect 179 280 181 285
rect 203 289 228 291
rect 203 281 205 289
rect 216 281 218 285
rect 226 281 228 289
rect 236 284 238 289
rect 243 284 245 289
rect 111 269 113 272
rect 104 267 113 269
rect 121 268 123 272
rect 131 269 133 272
rect 95 259 97 267
rect 104 265 106 267
rect 108 265 113 267
rect 104 263 113 265
rect 129 267 133 269
rect 129 264 131 267
rect 111 259 113 263
rect 125 262 131 264
rect 138 263 140 272
rect 200 279 205 281
rect 200 276 202 279
rect 159 264 161 269
rect 172 264 174 269
rect 125 260 127 262
rect 129 260 131 262
rect 92 257 105 259
rect 111 257 121 259
rect 125 258 131 260
rect 92 256 94 257
rect 74 254 80 256
rect 74 252 76 254
rect 78 252 80 254
rect 74 250 80 252
rect 88 254 94 256
rect 103 254 105 257
rect 119 254 121 257
rect 129 254 131 258
rect 135 261 141 263
rect 135 259 137 261
rect 139 259 141 261
rect 135 257 141 259
rect 139 254 141 257
rect 159 262 165 264
rect 159 260 161 262
rect 163 260 165 262
rect 159 258 165 260
rect 169 262 175 264
rect 169 260 171 262
rect 173 260 175 262
rect 169 258 175 260
rect 159 254 161 258
rect 88 252 90 254
rect 92 252 94 254
rect 88 250 94 252
rect 74 247 76 250
rect 54 232 56 236
rect 64 229 66 234
rect 74 229 76 234
rect 27 223 29 227
rect 34 223 36 227
rect 119 232 121 236
rect 129 232 131 236
rect 103 223 105 227
rect 169 247 171 258
rect 179 256 181 269
rect 216 269 218 272
rect 209 267 218 269
rect 226 268 228 272
rect 236 269 238 272
rect 200 259 202 267
rect 209 265 211 267
rect 213 265 218 267
rect 209 263 218 265
rect 234 267 238 269
rect 234 264 236 267
rect 216 259 218 263
rect 230 262 236 264
rect 243 263 245 272
rect 230 260 232 262
rect 234 260 236 262
rect 197 257 210 259
rect 216 257 226 259
rect 230 258 236 260
rect 197 256 199 257
rect 179 254 185 256
rect 179 252 181 254
rect 183 252 185 254
rect 179 250 185 252
rect 193 254 199 256
rect 208 254 210 257
rect 224 254 226 257
rect 234 254 236 258
rect 240 261 246 263
rect 240 259 242 261
rect 244 259 246 261
rect 240 257 246 259
rect 244 254 246 257
rect 193 252 195 254
rect 197 252 199 254
rect 193 250 199 252
rect 179 247 181 250
rect 159 232 161 236
rect 169 229 171 234
rect 179 229 181 234
rect 139 223 141 227
rect 224 232 226 236
rect 234 232 236 236
rect 208 223 210 227
rect 244 223 246 227
rect 27 215 29 219
rect 34 215 36 219
rect 14 205 16 210
rect 103 215 105 219
rect 54 206 56 210
rect 64 208 66 213
rect 74 208 76 213
rect 14 184 16 187
rect 27 184 29 194
rect 34 191 36 194
rect 34 189 40 191
rect 34 187 36 189
rect 38 187 40 189
rect 34 185 40 187
rect 14 182 20 184
rect 14 180 16 182
rect 18 180 20 182
rect 14 178 20 180
rect 24 182 30 184
rect 24 180 26 182
rect 28 180 30 182
rect 24 178 30 180
rect 14 175 16 178
rect 24 175 26 178
rect 34 175 36 185
rect 54 184 56 188
rect 64 184 66 195
rect 74 192 76 195
rect 74 190 80 192
rect 74 188 76 190
rect 78 188 80 190
rect 74 186 80 188
rect 88 190 94 192
rect 88 188 90 190
rect 92 188 94 190
rect 139 215 141 219
rect 119 206 121 210
rect 129 206 131 210
rect 208 215 210 219
rect 159 206 161 210
rect 169 208 171 213
rect 179 208 181 213
rect 88 186 94 188
rect 54 182 60 184
rect 54 180 56 182
rect 58 180 60 182
rect 54 178 60 180
rect 64 182 70 184
rect 64 180 66 182
rect 68 180 70 182
rect 64 178 70 180
rect 54 173 56 178
rect 67 173 69 178
rect 74 173 76 186
rect 92 185 94 186
rect 103 185 105 188
rect 119 185 121 188
rect 92 183 105 185
rect 111 183 121 185
rect 129 184 131 188
rect 139 185 141 188
rect 95 175 97 183
rect 111 179 113 183
rect 104 177 113 179
rect 125 182 131 184
rect 125 180 127 182
rect 129 180 131 182
rect 125 178 131 180
rect 135 183 141 185
rect 135 181 137 183
rect 139 181 141 183
rect 135 179 141 181
rect 159 184 161 188
rect 169 184 171 195
rect 179 192 181 195
rect 179 190 185 192
rect 179 188 181 190
rect 183 188 185 190
rect 179 186 185 188
rect 193 190 199 192
rect 193 188 195 190
rect 197 188 199 190
rect 244 215 246 219
rect 224 206 226 210
rect 234 206 236 210
rect 193 186 199 188
rect 159 182 165 184
rect 159 180 161 182
rect 163 180 165 182
rect 104 175 106 177
rect 108 175 113 177
rect 14 161 16 166
rect 24 164 26 169
rect 34 164 36 169
rect 54 160 56 164
rect 104 173 113 175
rect 129 175 131 178
rect 111 170 113 173
rect 121 170 123 174
rect 129 173 133 175
rect 131 170 133 173
rect 138 170 140 179
rect 159 178 165 180
rect 169 182 175 184
rect 169 180 171 182
rect 173 180 175 182
rect 169 178 175 180
rect 159 173 161 178
rect 172 173 174 178
rect 179 173 181 186
rect 197 185 199 186
rect 208 185 210 188
rect 224 185 226 188
rect 197 183 210 185
rect 216 183 226 185
rect 234 184 236 188
rect 244 185 246 188
rect 200 175 202 183
rect 216 179 218 183
rect 209 177 218 179
rect 230 182 236 184
rect 230 180 232 182
rect 234 180 236 182
rect 230 178 236 180
rect 240 183 246 185
rect 240 181 242 183
rect 244 181 246 183
rect 240 179 246 181
rect 209 175 211 177
rect 213 175 218 177
rect 95 163 97 166
rect 67 157 69 162
rect 74 157 76 162
rect 95 161 100 163
rect 98 153 100 161
rect 111 157 113 161
rect 121 153 123 161
rect 159 160 161 164
rect 209 173 218 175
rect 234 175 236 178
rect 216 170 218 173
rect 226 170 228 174
rect 234 173 238 175
rect 236 170 238 173
rect 243 170 245 179
rect 200 163 202 166
rect 131 153 133 158
rect 138 153 140 158
rect 98 151 123 153
rect 172 157 174 162
rect 179 157 181 162
rect 200 161 205 163
rect 203 153 205 161
rect 216 157 218 161
rect 226 153 228 161
rect 236 153 238 158
rect 243 153 245 158
rect 203 151 228 153
rect 14 132 16 137
rect 24 129 26 134
rect 34 129 36 134
rect 54 134 56 138
rect 67 136 69 141
rect 74 136 76 141
rect 98 145 123 147
rect 98 137 100 145
rect 111 137 113 141
rect 121 137 123 145
rect 131 140 133 145
rect 138 140 140 145
rect 95 135 100 137
rect 95 132 97 135
rect 14 120 16 123
rect 24 120 26 123
rect 14 118 20 120
rect 14 116 16 118
rect 18 116 20 118
rect 14 114 20 116
rect 24 118 30 120
rect 24 116 26 118
rect 28 116 30 118
rect 24 114 30 116
rect 14 111 16 114
rect 27 104 29 114
rect 34 113 36 123
rect 54 120 56 125
rect 67 120 69 125
rect 54 118 60 120
rect 54 116 56 118
rect 58 116 60 118
rect 54 114 60 116
rect 64 118 70 120
rect 64 116 66 118
rect 68 116 70 118
rect 64 114 70 116
rect 34 111 40 113
rect 34 109 36 111
rect 38 109 40 111
rect 54 110 56 114
rect 34 107 40 109
rect 34 104 36 107
rect 14 88 16 93
rect 64 103 66 114
rect 74 112 76 125
rect 159 134 161 138
rect 172 136 174 141
rect 179 136 181 141
rect 203 145 228 147
rect 203 137 205 145
rect 216 137 218 141
rect 226 137 228 145
rect 236 140 238 145
rect 243 140 245 145
rect 111 125 113 128
rect 104 123 113 125
rect 121 124 123 128
rect 131 125 133 128
rect 95 115 97 123
rect 104 121 106 123
rect 108 121 113 123
rect 104 119 113 121
rect 129 123 133 125
rect 129 120 131 123
rect 111 115 113 119
rect 125 118 131 120
rect 138 119 140 128
rect 200 135 205 137
rect 200 132 202 135
rect 159 120 161 125
rect 172 120 174 125
rect 125 116 127 118
rect 129 116 131 118
rect 92 113 105 115
rect 111 113 121 115
rect 125 114 131 116
rect 92 112 94 113
rect 74 110 80 112
rect 74 108 76 110
rect 78 108 80 110
rect 74 106 80 108
rect 88 110 94 112
rect 103 110 105 113
rect 119 110 121 113
rect 129 110 131 114
rect 135 117 141 119
rect 135 115 137 117
rect 139 115 141 117
rect 135 113 141 115
rect 139 110 141 113
rect 159 118 165 120
rect 159 116 161 118
rect 163 116 165 118
rect 159 114 165 116
rect 169 118 175 120
rect 169 116 171 118
rect 173 116 175 118
rect 169 114 175 116
rect 159 110 161 114
rect 88 108 90 110
rect 92 108 94 110
rect 88 106 94 108
rect 74 103 76 106
rect 54 88 56 92
rect 64 85 66 90
rect 74 85 76 90
rect 27 79 29 83
rect 34 79 36 83
rect 119 88 121 92
rect 129 88 131 92
rect 103 79 105 83
rect 169 103 171 114
rect 179 112 181 125
rect 216 125 218 128
rect 209 123 218 125
rect 226 124 228 128
rect 236 125 238 128
rect 200 115 202 123
rect 209 121 211 123
rect 213 121 218 123
rect 209 119 218 121
rect 234 123 238 125
rect 234 120 236 123
rect 216 115 218 119
rect 230 118 236 120
rect 243 119 245 128
rect 230 116 232 118
rect 234 116 236 118
rect 197 113 210 115
rect 216 113 226 115
rect 230 114 236 116
rect 197 112 199 113
rect 179 110 185 112
rect 179 108 181 110
rect 183 108 185 110
rect 179 106 185 108
rect 193 110 199 112
rect 208 110 210 113
rect 224 110 226 113
rect 234 110 236 114
rect 240 117 246 119
rect 240 115 242 117
rect 244 115 246 117
rect 240 113 246 115
rect 244 110 246 113
rect 193 108 195 110
rect 197 108 199 110
rect 193 106 199 108
rect 179 103 181 106
rect 159 88 161 92
rect 169 85 171 90
rect 179 85 181 90
rect 139 79 141 83
rect 224 88 226 92
rect 234 88 236 92
rect 208 79 210 83
rect 244 79 246 83
rect 27 71 29 75
rect 34 71 36 75
rect 14 61 16 66
rect 103 71 105 75
rect 54 62 56 66
rect 64 64 66 69
rect 74 64 76 69
rect 14 40 16 43
rect 27 40 29 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 31 16 34
rect 24 31 26 34
rect 34 31 36 41
rect 54 40 56 44
rect 64 40 66 51
rect 74 48 76 51
rect 74 46 80 48
rect 74 44 76 46
rect 78 44 80 46
rect 74 42 80 44
rect 88 46 94 48
rect 88 44 90 46
rect 92 44 94 46
rect 139 71 141 75
rect 119 62 121 66
rect 129 62 131 66
rect 208 71 210 75
rect 159 62 161 66
rect 169 64 171 69
rect 179 64 181 69
rect 88 42 94 44
rect 54 38 60 40
rect 54 36 56 38
rect 58 36 60 38
rect 54 34 60 36
rect 64 38 70 40
rect 64 36 66 38
rect 68 36 70 38
rect 64 34 70 36
rect 54 29 56 34
rect 67 29 69 34
rect 74 29 76 42
rect 92 41 94 42
rect 103 41 105 44
rect 119 41 121 44
rect 92 39 105 41
rect 111 39 121 41
rect 129 40 131 44
rect 139 41 141 44
rect 95 31 97 39
rect 111 35 113 39
rect 104 33 113 35
rect 125 38 131 40
rect 125 36 127 38
rect 129 36 131 38
rect 125 34 131 36
rect 135 39 141 41
rect 135 37 137 39
rect 139 37 141 39
rect 135 35 141 37
rect 159 40 161 44
rect 169 40 171 51
rect 179 48 181 51
rect 179 46 185 48
rect 179 44 181 46
rect 183 44 185 46
rect 179 42 185 44
rect 193 46 199 48
rect 193 44 195 46
rect 197 44 199 46
rect 244 71 246 75
rect 224 62 226 66
rect 234 62 236 66
rect 193 42 199 44
rect 159 38 165 40
rect 159 36 161 38
rect 163 36 165 38
rect 104 31 106 33
rect 108 31 113 33
rect 14 17 16 22
rect 24 20 26 25
rect 34 20 36 25
rect 54 16 56 20
rect 104 29 113 31
rect 129 31 131 34
rect 111 26 113 29
rect 121 26 123 30
rect 129 29 133 31
rect 131 26 133 29
rect 138 26 140 35
rect 159 34 165 36
rect 169 38 175 40
rect 169 36 171 38
rect 173 36 175 38
rect 169 34 175 36
rect 159 29 161 34
rect 172 29 174 34
rect 179 29 181 42
rect 197 41 199 42
rect 208 41 210 44
rect 224 41 226 44
rect 197 39 210 41
rect 216 39 226 41
rect 234 40 236 44
rect 244 41 246 44
rect 200 31 202 39
rect 216 35 218 39
rect 209 33 218 35
rect 230 38 236 40
rect 230 36 232 38
rect 234 36 236 38
rect 230 34 236 36
rect 240 39 246 41
rect 240 37 242 39
rect 244 37 246 39
rect 240 35 246 37
rect 209 31 211 33
rect 213 31 218 33
rect 95 19 97 22
rect 67 13 69 18
rect 74 13 76 18
rect 95 17 100 19
rect 98 9 100 17
rect 111 13 113 17
rect 121 9 123 17
rect 159 16 161 20
rect 209 29 218 31
rect 234 31 236 34
rect 216 26 218 29
rect 226 26 228 30
rect 234 29 238 31
rect 236 26 238 29
rect 243 26 245 35
rect 200 19 202 22
rect 131 9 133 14
rect 138 9 140 14
rect 98 7 123 9
rect 172 13 174 18
rect 179 13 181 18
rect 200 17 205 19
rect 203 9 205 17
rect 216 13 218 17
rect 226 9 228 17
rect 236 9 238 14
rect 243 9 245 14
rect 203 7 228 9
<< ndif >>
rect 18 284 24 286
rect 18 282 20 284
rect 22 282 24 284
rect 18 280 24 282
rect 37 284 43 286
rect 58 288 65 290
rect 58 286 60 288
rect 62 286 65 288
rect 37 282 39 284
rect 41 282 43 284
rect 37 280 43 282
rect 18 276 22 280
rect 9 273 14 276
rect 7 271 14 273
rect 7 269 9 271
rect 11 269 14 271
rect 7 267 14 269
rect 16 273 22 276
rect 38 273 43 280
rect 58 280 65 286
rect 142 288 148 290
rect 142 286 144 288
rect 146 286 148 288
rect 142 284 148 286
rect 163 288 170 290
rect 163 286 165 288
rect 167 286 170 288
rect 126 281 131 284
rect 58 278 67 280
rect 16 267 24 273
rect 26 271 34 273
rect 26 269 29 271
rect 31 269 34 271
rect 26 267 34 269
rect 36 267 43 273
rect 47 276 54 278
rect 47 274 49 276
rect 51 274 54 276
rect 47 272 54 274
rect 49 269 54 272
rect 56 269 67 278
rect 69 269 74 280
rect 76 278 83 280
rect 76 276 79 278
rect 81 276 83 278
rect 102 279 111 281
rect 102 277 104 279
rect 106 277 111 279
rect 102 276 111 277
rect 76 274 83 276
rect 76 269 81 274
rect 90 273 95 276
rect 88 271 95 273
rect 88 269 90 271
rect 92 269 95 271
rect 88 267 95 269
rect 97 272 111 276
rect 113 276 121 281
rect 113 274 116 276
rect 118 274 121 276
rect 113 272 121 274
rect 123 278 131 281
rect 123 276 126 278
rect 128 276 131 278
rect 123 272 131 276
rect 133 272 138 284
rect 140 272 148 284
rect 163 280 170 286
rect 247 288 253 290
rect 247 286 249 288
rect 251 286 253 288
rect 247 284 253 286
rect 231 281 236 284
rect 163 278 172 280
rect 152 276 159 278
rect 152 274 154 276
rect 156 274 159 276
rect 152 272 159 274
rect 97 267 102 272
rect 154 269 159 272
rect 161 269 172 278
rect 174 269 179 280
rect 181 278 188 280
rect 181 276 184 278
rect 186 276 188 278
rect 207 279 216 281
rect 207 277 209 279
rect 211 277 216 279
rect 207 276 216 277
rect 181 274 188 276
rect 181 269 186 274
rect 195 273 200 276
rect 193 271 200 273
rect 193 269 195 271
rect 197 269 200 271
rect 193 267 200 269
rect 202 272 216 276
rect 218 276 226 281
rect 218 274 221 276
rect 223 274 226 276
rect 218 272 226 274
rect 228 278 236 281
rect 228 276 231 278
rect 233 276 236 278
rect 228 272 236 276
rect 238 272 243 284
rect 245 272 253 284
rect 202 267 207 272
rect 7 173 14 175
rect 7 171 9 173
rect 11 171 14 173
rect 7 169 14 171
rect 9 166 14 169
rect 16 169 24 175
rect 26 173 34 175
rect 26 171 29 173
rect 31 171 34 173
rect 26 169 34 171
rect 36 169 43 175
rect 88 173 95 175
rect 49 170 54 173
rect 16 166 22 169
rect 18 162 22 166
rect 38 162 43 169
rect 47 168 54 170
rect 47 166 49 168
rect 51 166 54 168
rect 47 164 54 166
rect 56 164 67 173
rect 18 160 24 162
rect 18 158 20 160
rect 22 158 24 160
rect 18 156 24 158
rect 37 160 43 162
rect 58 162 67 164
rect 69 162 74 173
rect 76 168 81 173
rect 88 171 90 173
rect 92 171 95 173
rect 88 169 95 171
rect 76 166 83 168
rect 90 166 95 169
rect 97 170 102 175
rect 193 173 200 175
rect 154 170 159 173
rect 97 166 111 170
rect 76 164 79 166
rect 81 164 83 166
rect 76 162 83 164
rect 102 165 111 166
rect 102 163 104 165
rect 106 163 111 165
rect 37 158 39 160
rect 41 158 43 160
rect 37 156 43 158
rect 58 156 65 162
rect 102 161 111 163
rect 113 168 121 170
rect 113 166 116 168
rect 118 166 121 168
rect 113 161 121 166
rect 123 166 131 170
rect 123 164 126 166
rect 128 164 131 166
rect 123 161 131 164
rect 58 154 60 156
rect 62 154 65 156
rect 58 152 65 154
rect 126 158 131 161
rect 133 158 138 170
rect 140 158 148 170
rect 152 168 159 170
rect 152 166 154 168
rect 156 166 159 168
rect 152 164 159 166
rect 161 164 172 173
rect 163 162 172 164
rect 174 162 179 173
rect 181 168 186 173
rect 193 171 195 173
rect 197 171 200 173
rect 193 169 200 171
rect 181 166 188 168
rect 195 166 200 169
rect 202 170 207 175
rect 202 166 216 170
rect 181 164 184 166
rect 186 164 188 166
rect 181 162 188 164
rect 207 165 216 166
rect 207 163 209 165
rect 211 163 216 165
rect 142 156 148 158
rect 142 154 144 156
rect 146 154 148 156
rect 142 152 148 154
rect 163 156 170 162
rect 207 161 216 163
rect 218 168 226 170
rect 218 166 221 168
rect 223 166 226 168
rect 218 161 226 166
rect 228 166 236 170
rect 228 164 231 166
rect 233 164 236 166
rect 228 161 236 164
rect 163 154 165 156
rect 167 154 170 156
rect 163 152 170 154
rect 231 158 236 161
rect 238 158 243 170
rect 245 158 253 170
rect 247 156 253 158
rect 247 154 249 156
rect 251 154 253 156
rect 247 152 253 154
rect 18 140 24 142
rect 18 138 20 140
rect 22 138 24 140
rect 18 136 24 138
rect 37 140 43 142
rect 58 144 65 146
rect 58 142 60 144
rect 62 142 65 144
rect 37 138 39 140
rect 41 138 43 140
rect 37 136 43 138
rect 18 132 22 136
rect 9 129 14 132
rect 7 127 14 129
rect 7 125 9 127
rect 11 125 14 127
rect 7 123 14 125
rect 16 129 22 132
rect 38 129 43 136
rect 58 136 65 142
rect 142 144 148 146
rect 142 142 144 144
rect 146 142 148 144
rect 142 140 148 142
rect 163 144 170 146
rect 163 142 165 144
rect 167 142 170 144
rect 126 137 131 140
rect 58 134 67 136
rect 16 123 24 129
rect 26 127 34 129
rect 26 125 29 127
rect 31 125 34 127
rect 26 123 34 125
rect 36 123 43 129
rect 47 132 54 134
rect 47 130 49 132
rect 51 130 54 132
rect 47 128 54 130
rect 49 125 54 128
rect 56 125 67 134
rect 69 125 74 136
rect 76 134 83 136
rect 76 132 79 134
rect 81 132 83 134
rect 102 135 111 137
rect 102 133 104 135
rect 106 133 111 135
rect 102 132 111 133
rect 76 130 83 132
rect 76 125 81 130
rect 90 129 95 132
rect 88 127 95 129
rect 88 125 90 127
rect 92 125 95 127
rect 88 123 95 125
rect 97 128 111 132
rect 113 132 121 137
rect 113 130 116 132
rect 118 130 121 132
rect 113 128 121 130
rect 123 134 131 137
rect 123 132 126 134
rect 128 132 131 134
rect 123 128 131 132
rect 133 128 138 140
rect 140 128 148 140
rect 163 136 170 142
rect 247 144 253 146
rect 247 142 249 144
rect 251 142 253 144
rect 247 140 253 142
rect 231 137 236 140
rect 163 134 172 136
rect 152 132 159 134
rect 152 130 154 132
rect 156 130 159 132
rect 152 128 159 130
rect 97 123 102 128
rect 154 125 159 128
rect 161 125 172 134
rect 174 125 179 136
rect 181 134 188 136
rect 181 132 184 134
rect 186 132 188 134
rect 207 135 216 137
rect 207 133 209 135
rect 211 133 216 135
rect 207 132 216 133
rect 181 130 188 132
rect 181 125 186 130
rect 195 129 200 132
rect 193 127 200 129
rect 193 125 195 127
rect 197 125 200 127
rect 193 123 200 125
rect 202 128 216 132
rect 218 132 226 137
rect 218 130 221 132
rect 223 130 226 132
rect 218 128 226 130
rect 228 134 236 137
rect 228 132 231 134
rect 233 132 236 134
rect 228 128 236 132
rect 238 128 243 140
rect 245 128 253 140
rect 202 123 207 128
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 9 22 14 25
rect 16 25 24 31
rect 26 29 34 31
rect 26 27 29 29
rect 31 27 34 29
rect 26 25 34 27
rect 36 25 43 31
rect 88 29 95 31
rect 49 26 54 29
rect 16 22 22 25
rect 18 18 22 22
rect 38 18 43 25
rect 47 24 54 26
rect 47 22 49 24
rect 51 22 54 24
rect 47 20 54 22
rect 56 20 67 29
rect 18 16 24 18
rect 18 14 20 16
rect 22 14 24 16
rect 18 12 24 14
rect 37 16 43 18
rect 58 18 67 20
rect 69 18 74 29
rect 76 24 81 29
rect 88 27 90 29
rect 92 27 95 29
rect 88 25 95 27
rect 76 22 83 24
rect 90 22 95 25
rect 97 26 102 31
rect 193 29 200 31
rect 154 26 159 29
rect 97 22 111 26
rect 76 20 79 22
rect 81 20 83 22
rect 76 18 83 20
rect 102 21 111 22
rect 102 19 104 21
rect 106 19 111 21
rect 37 14 39 16
rect 41 14 43 16
rect 37 12 43 14
rect 58 12 65 18
rect 102 17 111 19
rect 113 24 121 26
rect 113 22 116 24
rect 118 22 121 24
rect 113 17 121 22
rect 123 22 131 26
rect 123 20 126 22
rect 128 20 131 22
rect 123 17 131 20
rect 58 10 60 12
rect 62 10 65 12
rect 58 8 65 10
rect 126 14 131 17
rect 133 14 138 26
rect 140 14 148 26
rect 152 24 159 26
rect 152 22 154 24
rect 156 22 159 24
rect 152 20 159 22
rect 161 20 172 29
rect 163 18 172 20
rect 174 18 179 29
rect 181 24 186 29
rect 193 27 195 29
rect 197 27 200 29
rect 193 25 200 27
rect 181 22 188 24
rect 195 22 200 25
rect 202 26 207 31
rect 202 22 216 26
rect 181 20 184 22
rect 186 20 188 22
rect 181 18 188 20
rect 207 21 216 22
rect 207 19 209 21
rect 211 19 216 21
rect 142 12 148 14
rect 142 10 144 12
rect 146 10 148 12
rect 142 8 148 10
rect 163 12 170 18
rect 207 17 216 19
rect 218 24 226 26
rect 218 22 221 24
rect 223 22 226 24
rect 218 17 226 22
rect 228 22 236 26
rect 228 20 231 22
rect 233 20 236 22
rect 228 17 236 20
rect 163 10 165 12
rect 167 10 170 12
rect 163 8 170 10
rect 231 14 236 17
rect 238 14 243 26
rect 245 14 253 26
rect 247 12 253 14
rect 247 10 249 12
rect 251 10 253 12
rect 247 8 253 10
<< pdif >>
rect 9 250 14 255
rect 7 248 14 250
rect 7 246 9 248
rect 11 246 14 248
rect 7 241 14 246
rect 7 239 9 241
rect 11 239 14 241
rect 7 237 14 239
rect 16 248 24 255
rect 47 252 54 254
rect 47 250 49 252
rect 51 250 54 252
rect 16 237 27 248
rect 18 231 27 237
rect 18 229 20 231
rect 22 229 27 231
rect 18 227 27 229
rect 29 227 34 248
rect 36 240 41 248
rect 47 245 54 250
rect 47 243 49 245
rect 51 243 54 245
rect 47 241 54 243
rect 36 238 43 240
rect 36 236 39 238
rect 41 236 43 238
rect 49 236 54 241
rect 56 247 62 254
rect 96 252 103 254
rect 96 250 98 252
rect 100 250 103 252
rect 96 248 103 250
rect 56 240 64 247
rect 56 238 59 240
rect 61 238 64 240
rect 56 236 64 238
rect 36 234 43 236
rect 36 227 41 234
rect 58 234 64 236
rect 66 245 74 247
rect 66 243 69 245
rect 71 243 74 245
rect 66 238 74 243
rect 66 236 69 238
rect 71 236 74 238
rect 66 234 74 236
rect 76 238 83 247
rect 76 236 79 238
rect 81 236 83 238
rect 76 234 83 236
rect 98 227 103 248
rect 105 238 119 254
rect 105 236 108 238
rect 110 236 119 238
rect 121 252 129 254
rect 121 250 124 252
rect 126 250 129 252
rect 121 245 129 250
rect 121 243 124 245
rect 126 243 129 245
rect 121 236 129 243
rect 131 245 139 254
rect 131 243 134 245
rect 136 243 139 245
rect 131 236 139 243
rect 105 231 117 236
rect 105 229 108 231
rect 110 229 117 231
rect 105 227 117 229
rect 134 227 139 236
rect 141 239 146 254
rect 152 252 159 254
rect 152 250 154 252
rect 156 250 159 252
rect 152 245 159 250
rect 152 243 154 245
rect 156 243 159 245
rect 152 241 159 243
rect 141 237 148 239
rect 141 235 144 237
rect 146 235 148 237
rect 154 236 159 241
rect 161 247 167 254
rect 201 252 208 254
rect 201 250 203 252
rect 205 250 208 252
rect 201 248 208 250
rect 161 240 169 247
rect 161 238 164 240
rect 166 238 169 240
rect 161 236 169 238
rect 141 233 148 235
rect 141 227 146 233
rect 163 234 169 236
rect 171 245 179 247
rect 171 243 174 245
rect 176 243 179 245
rect 171 238 179 243
rect 171 236 174 238
rect 176 236 179 238
rect 171 234 179 236
rect 181 238 188 247
rect 181 236 184 238
rect 186 236 188 238
rect 181 234 188 236
rect 203 227 208 248
rect 210 238 224 254
rect 210 236 213 238
rect 215 236 224 238
rect 226 252 234 254
rect 226 250 229 252
rect 231 250 234 252
rect 226 245 234 250
rect 226 243 229 245
rect 231 243 234 245
rect 226 236 234 243
rect 236 245 244 254
rect 236 243 239 245
rect 241 243 244 245
rect 236 236 244 243
rect 210 231 222 236
rect 210 229 213 231
rect 215 229 222 231
rect 210 227 222 229
rect 239 227 244 236
rect 246 239 251 254
rect 246 237 253 239
rect 246 235 249 237
rect 251 235 253 237
rect 246 233 253 235
rect 246 227 251 233
rect 18 213 27 215
rect 18 211 20 213
rect 22 211 27 213
rect 18 205 27 211
rect 7 203 14 205
rect 7 201 9 203
rect 11 201 14 203
rect 7 196 14 201
rect 7 194 9 196
rect 11 194 14 196
rect 7 192 14 194
rect 9 187 14 192
rect 16 194 27 205
rect 29 194 34 215
rect 36 208 41 215
rect 36 206 43 208
rect 58 206 64 208
rect 36 204 39 206
rect 41 204 43 206
rect 36 202 43 204
rect 36 194 41 202
rect 49 201 54 206
rect 47 199 54 201
rect 47 197 49 199
rect 51 197 54 199
rect 16 187 24 194
rect 47 192 54 197
rect 47 190 49 192
rect 51 190 54 192
rect 47 188 54 190
rect 56 204 64 206
rect 56 202 59 204
rect 61 202 64 204
rect 56 195 64 202
rect 66 206 74 208
rect 66 204 69 206
rect 71 204 74 206
rect 66 199 74 204
rect 66 197 69 199
rect 71 197 74 199
rect 66 195 74 197
rect 76 206 83 208
rect 76 204 79 206
rect 81 204 83 206
rect 76 195 83 204
rect 56 188 62 195
rect 98 194 103 215
rect 96 192 103 194
rect 96 190 98 192
rect 100 190 103 192
rect 96 188 103 190
rect 105 213 117 215
rect 105 211 108 213
rect 110 211 117 213
rect 105 206 117 211
rect 134 206 139 215
rect 105 204 108 206
rect 110 204 119 206
rect 105 188 119 204
rect 121 199 129 206
rect 121 197 124 199
rect 126 197 129 199
rect 121 192 129 197
rect 121 190 124 192
rect 126 190 129 192
rect 121 188 129 190
rect 131 199 139 206
rect 131 197 134 199
rect 136 197 139 199
rect 131 188 139 197
rect 141 209 146 215
rect 141 207 148 209
rect 141 205 144 207
rect 146 205 148 207
rect 163 206 169 208
rect 141 203 148 205
rect 141 188 146 203
rect 154 201 159 206
rect 152 199 159 201
rect 152 197 154 199
rect 156 197 159 199
rect 152 192 159 197
rect 152 190 154 192
rect 156 190 159 192
rect 152 188 159 190
rect 161 204 169 206
rect 161 202 164 204
rect 166 202 169 204
rect 161 195 169 202
rect 171 206 179 208
rect 171 204 174 206
rect 176 204 179 206
rect 171 199 179 204
rect 171 197 174 199
rect 176 197 179 199
rect 171 195 179 197
rect 181 206 188 208
rect 181 204 184 206
rect 186 204 188 206
rect 181 195 188 204
rect 161 188 167 195
rect 203 194 208 215
rect 201 192 208 194
rect 201 190 203 192
rect 205 190 208 192
rect 201 188 208 190
rect 210 213 222 215
rect 210 211 213 213
rect 215 211 222 213
rect 210 206 222 211
rect 239 206 244 215
rect 210 204 213 206
rect 215 204 224 206
rect 210 188 224 204
rect 226 199 234 206
rect 226 197 229 199
rect 231 197 234 199
rect 226 192 234 197
rect 226 190 229 192
rect 231 190 234 192
rect 226 188 234 190
rect 236 199 244 206
rect 236 197 239 199
rect 241 197 244 199
rect 236 188 244 197
rect 246 209 251 215
rect 246 207 253 209
rect 246 205 249 207
rect 251 205 253 207
rect 246 203 253 205
rect 246 188 251 203
rect 9 106 14 111
rect 7 104 14 106
rect 7 102 9 104
rect 11 102 14 104
rect 7 97 14 102
rect 7 95 9 97
rect 11 95 14 97
rect 7 93 14 95
rect 16 104 24 111
rect 47 108 54 110
rect 47 106 49 108
rect 51 106 54 108
rect 16 93 27 104
rect 18 87 27 93
rect 18 85 20 87
rect 22 85 27 87
rect 18 83 27 85
rect 29 83 34 104
rect 36 96 41 104
rect 47 101 54 106
rect 47 99 49 101
rect 51 99 54 101
rect 47 97 54 99
rect 36 94 43 96
rect 36 92 39 94
rect 41 92 43 94
rect 49 92 54 97
rect 56 103 62 110
rect 96 108 103 110
rect 96 106 98 108
rect 100 106 103 108
rect 96 104 103 106
rect 56 96 64 103
rect 56 94 59 96
rect 61 94 64 96
rect 56 92 64 94
rect 36 90 43 92
rect 36 83 41 90
rect 58 90 64 92
rect 66 101 74 103
rect 66 99 69 101
rect 71 99 74 101
rect 66 94 74 99
rect 66 92 69 94
rect 71 92 74 94
rect 66 90 74 92
rect 76 94 83 103
rect 76 92 79 94
rect 81 92 83 94
rect 76 90 83 92
rect 98 83 103 104
rect 105 94 119 110
rect 105 92 108 94
rect 110 92 119 94
rect 121 108 129 110
rect 121 106 124 108
rect 126 106 129 108
rect 121 101 129 106
rect 121 99 124 101
rect 126 99 129 101
rect 121 92 129 99
rect 131 101 139 110
rect 131 99 134 101
rect 136 99 139 101
rect 131 92 139 99
rect 105 87 117 92
rect 105 85 108 87
rect 110 85 117 87
rect 105 83 117 85
rect 134 83 139 92
rect 141 95 146 110
rect 152 108 159 110
rect 152 106 154 108
rect 156 106 159 108
rect 152 101 159 106
rect 152 99 154 101
rect 156 99 159 101
rect 152 97 159 99
rect 141 93 148 95
rect 141 91 144 93
rect 146 91 148 93
rect 154 92 159 97
rect 161 103 167 110
rect 201 108 208 110
rect 201 106 203 108
rect 205 106 208 108
rect 201 104 208 106
rect 161 96 169 103
rect 161 94 164 96
rect 166 94 169 96
rect 161 92 169 94
rect 141 89 148 91
rect 141 83 146 89
rect 163 90 169 92
rect 171 101 179 103
rect 171 99 174 101
rect 176 99 179 101
rect 171 94 179 99
rect 171 92 174 94
rect 176 92 179 94
rect 171 90 179 92
rect 181 94 188 103
rect 181 92 184 94
rect 186 92 188 94
rect 181 90 188 92
rect 203 83 208 104
rect 210 94 224 110
rect 210 92 213 94
rect 215 92 224 94
rect 226 108 234 110
rect 226 106 229 108
rect 231 106 234 108
rect 226 101 234 106
rect 226 99 229 101
rect 231 99 234 101
rect 226 92 234 99
rect 236 101 244 110
rect 236 99 239 101
rect 241 99 244 101
rect 236 92 244 99
rect 210 87 222 92
rect 210 85 213 87
rect 215 85 222 87
rect 210 83 222 85
rect 239 83 244 92
rect 246 95 251 110
rect 246 93 253 95
rect 246 91 249 93
rect 251 91 253 93
rect 246 89 253 91
rect 246 83 251 89
rect 18 69 27 71
rect 18 67 20 69
rect 22 67 27 69
rect 18 61 27 67
rect 7 59 14 61
rect 7 57 9 59
rect 11 57 14 59
rect 7 52 14 57
rect 7 50 9 52
rect 11 50 14 52
rect 7 48 14 50
rect 9 43 14 48
rect 16 50 27 61
rect 29 50 34 71
rect 36 64 41 71
rect 36 62 43 64
rect 58 62 64 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 58 43 60
rect 36 50 41 58
rect 49 57 54 62
rect 47 55 54 57
rect 47 53 49 55
rect 51 53 54 55
rect 16 43 24 50
rect 47 48 54 53
rect 47 46 49 48
rect 51 46 54 48
rect 47 44 54 46
rect 56 60 64 62
rect 56 58 59 60
rect 61 58 64 60
rect 56 51 64 58
rect 66 62 74 64
rect 66 60 69 62
rect 71 60 74 62
rect 66 55 74 60
rect 66 53 69 55
rect 71 53 74 55
rect 66 51 74 53
rect 76 62 83 64
rect 76 60 79 62
rect 81 60 83 62
rect 76 51 83 60
rect 56 44 62 51
rect 98 50 103 71
rect 96 48 103 50
rect 96 46 98 48
rect 100 46 103 48
rect 96 44 103 46
rect 105 69 117 71
rect 105 67 108 69
rect 110 67 117 69
rect 105 62 117 67
rect 134 62 139 71
rect 105 60 108 62
rect 110 60 119 62
rect 105 44 119 60
rect 121 55 129 62
rect 121 53 124 55
rect 126 53 129 55
rect 121 48 129 53
rect 121 46 124 48
rect 126 46 129 48
rect 121 44 129 46
rect 131 55 139 62
rect 131 53 134 55
rect 136 53 139 55
rect 131 44 139 53
rect 141 65 146 71
rect 141 63 148 65
rect 141 61 144 63
rect 146 61 148 63
rect 163 62 169 64
rect 141 59 148 61
rect 141 44 146 59
rect 154 57 159 62
rect 152 55 159 57
rect 152 53 154 55
rect 156 53 159 55
rect 152 48 159 53
rect 152 46 154 48
rect 156 46 159 48
rect 152 44 159 46
rect 161 60 169 62
rect 161 58 164 60
rect 166 58 169 60
rect 161 51 169 58
rect 171 62 179 64
rect 171 60 174 62
rect 176 60 179 62
rect 171 55 179 60
rect 171 53 174 55
rect 176 53 179 55
rect 171 51 179 53
rect 181 62 188 64
rect 181 60 184 62
rect 186 60 188 62
rect 181 51 188 60
rect 161 44 167 51
rect 203 50 208 71
rect 201 48 208 50
rect 201 46 203 48
rect 205 46 208 48
rect 201 44 208 46
rect 210 69 222 71
rect 210 67 213 69
rect 215 67 222 69
rect 210 62 222 67
rect 239 62 244 71
rect 210 60 213 62
rect 215 60 224 62
rect 210 44 224 60
rect 226 55 234 62
rect 226 53 229 55
rect 231 53 234 55
rect 226 48 234 53
rect 226 46 229 48
rect 231 46 234 48
rect 226 44 234 46
rect 236 55 244 62
rect 236 53 239 55
rect 241 53 244 55
rect 236 44 244 53
rect 246 65 251 71
rect 246 63 253 65
rect 246 61 249 63
rect 251 61 253 63
rect 246 59 253 61
rect 246 44 251 59
<< alu1 >>
rect 3 288 257 293
rect 3 286 10 288
rect 12 286 50 288
rect 52 286 60 288
rect 62 286 91 288
rect 93 286 144 288
rect 146 286 155 288
rect 157 286 165 288
rect 167 286 196 288
rect 198 286 249 288
rect 251 286 257 288
rect 3 285 257 286
rect 47 276 59 280
rect 47 274 49 276
rect 51 274 59 276
rect 124 278 148 279
rect 7 271 12 273
rect 7 269 9 271
rect 11 269 12 271
rect 7 267 12 269
rect 7 248 11 267
rect 39 263 43 272
rect 47 263 51 274
rect 124 276 126 278
rect 128 276 148 278
rect 124 275 148 276
rect 7 246 9 248
rect 7 241 11 246
rect 7 239 9 241
rect 22 262 51 263
rect 22 260 26 262
rect 28 260 51 262
rect 22 259 51 260
rect 22 253 36 255
rect 38 253 43 255
rect 22 251 43 253
rect 39 245 43 251
rect 39 243 40 245
rect 42 243 43 245
rect 39 242 43 243
rect 47 254 51 259
rect 71 271 76 272
rect 71 269 72 271
rect 74 269 76 271
rect 71 263 76 269
rect 47 252 52 254
rect 47 250 49 252
rect 51 250 52 252
rect 47 245 52 250
rect 47 243 49 245
rect 51 243 52 245
rect 62 262 76 263
rect 62 260 66 262
rect 68 260 76 262
rect 62 259 76 260
rect 96 271 109 272
rect 96 269 99 271
rect 101 269 109 271
rect 96 267 109 269
rect 144 271 148 275
rect 96 266 106 267
rect 104 265 106 266
rect 108 265 109 267
rect 88 255 93 256
rect 70 254 83 255
rect 87 254 93 255
rect 70 252 76 254
rect 78 252 90 254
rect 92 252 93 254
rect 70 251 93 252
rect 79 249 93 251
rect 104 258 109 265
rect 144 269 145 271
rect 147 269 148 271
rect 47 241 52 243
rect 7 235 20 239
rect 7 234 11 235
rect 79 242 83 249
rect 88 240 93 249
rect 88 234 100 240
rect 144 247 148 269
rect 132 245 148 247
rect 132 243 134 245
rect 136 243 148 245
rect 132 242 148 243
rect 152 276 164 280
rect 152 274 154 276
rect 156 274 164 276
rect 229 278 253 279
rect 152 254 156 274
rect 229 276 231 278
rect 233 276 253 278
rect 229 275 253 276
rect 176 271 181 272
rect 176 269 177 271
rect 179 269 181 271
rect 176 263 181 269
rect 152 252 157 254
rect 152 250 154 252
rect 156 250 157 252
rect 152 245 157 250
rect 152 243 154 245
rect 156 243 157 245
rect 167 262 181 263
rect 167 260 171 262
rect 173 260 181 262
rect 167 259 181 260
rect 201 271 214 272
rect 201 269 204 271
rect 206 269 214 271
rect 201 267 214 269
rect 201 266 211 267
rect 209 265 211 266
rect 213 265 214 267
rect 193 255 198 256
rect 175 254 188 255
rect 192 254 198 255
rect 175 252 181 254
rect 183 252 195 254
rect 197 252 198 254
rect 175 251 198 252
rect 184 249 198 251
rect 209 258 214 265
rect 152 241 157 243
rect 184 246 188 249
rect 184 244 185 246
rect 187 244 188 246
rect 184 242 188 244
rect 193 240 198 249
rect 193 234 205 240
rect 249 247 253 275
rect 237 245 253 247
rect 237 243 239 245
rect 241 243 253 245
rect 237 242 253 243
rect 3 228 257 229
rect 3 226 10 228
rect 12 226 50 228
rect 52 226 124 228
rect 126 226 155 228
rect 157 226 229 228
rect 231 226 257 228
rect 3 216 257 226
rect 3 214 10 216
rect 12 214 50 216
rect 52 214 124 216
rect 126 214 155 216
rect 157 214 229 216
rect 231 214 257 216
rect 3 213 257 214
rect 7 207 11 208
rect 7 205 8 207
rect 10 205 20 207
rect 7 203 20 205
rect 7 201 9 203
rect 7 196 11 201
rect 7 194 9 196
rect 7 175 11 194
rect 39 199 43 200
rect 39 197 40 199
rect 42 197 43 199
rect 39 191 43 197
rect 22 189 43 191
rect 22 187 36 189
rect 38 187 43 189
rect 47 199 52 201
rect 47 197 49 199
rect 51 197 52 199
rect 88 202 100 208
rect 47 192 52 197
rect 47 190 49 192
rect 51 190 52 192
rect 47 188 52 190
rect 47 183 51 188
rect 7 173 12 175
rect 7 171 9 173
rect 11 171 12 173
rect 7 169 12 171
rect 22 182 51 183
rect 22 180 26 182
rect 28 180 51 182
rect 22 179 51 180
rect 39 170 43 179
rect 47 168 51 179
rect 79 193 83 200
rect 88 193 93 202
rect 79 191 93 193
rect 70 190 93 191
rect 70 188 76 190
rect 78 188 90 190
rect 92 188 93 190
rect 70 187 83 188
rect 87 187 93 188
rect 88 186 93 187
rect 62 182 76 183
rect 62 180 66 182
rect 68 180 76 182
rect 62 179 76 180
rect 47 166 49 168
rect 51 166 59 168
rect 47 162 59 166
rect 71 173 76 179
rect 71 171 72 173
rect 74 171 76 173
rect 71 170 76 171
rect 104 177 109 184
rect 132 199 148 200
rect 132 197 134 199
rect 136 197 148 199
rect 132 195 148 197
rect 104 176 106 177
rect 96 175 106 176
rect 108 175 109 177
rect 96 173 109 175
rect 96 171 99 173
rect 101 171 109 173
rect 96 170 109 171
rect 144 173 148 195
rect 144 171 145 173
rect 147 171 148 173
rect 144 167 148 171
rect 124 166 148 167
rect 124 164 126 166
rect 128 164 148 166
rect 124 163 148 164
rect 152 199 157 201
rect 152 197 154 199
rect 156 197 157 199
rect 193 202 205 208
rect 152 192 157 197
rect 152 190 154 192
rect 156 190 157 192
rect 152 188 157 190
rect 152 168 156 188
rect 184 193 188 200
rect 193 193 198 202
rect 184 191 198 193
rect 175 190 198 191
rect 175 188 176 190
rect 178 188 181 190
rect 183 188 195 190
rect 197 188 198 190
rect 175 187 188 188
rect 192 187 198 188
rect 193 186 198 187
rect 167 182 181 183
rect 167 180 171 182
rect 173 180 181 182
rect 167 179 181 180
rect 152 166 154 168
rect 156 166 164 168
rect 152 162 164 166
rect 176 173 181 179
rect 176 171 177 173
rect 179 171 181 173
rect 176 170 181 171
rect 209 177 214 184
rect 237 199 253 200
rect 237 197 239 199
rect 241 197 253 199
rect 237 195 253 197
rect 209 176 211 177
rect 201 175 211 176
rect 213 175 214 177
rect 201 173 214 175
rect 201 171 204 173
rect 206 171 214 173
rect 201 170 214 171
rect 249 167 253 195
rect 229 166 253 167
rect 229 164 231 166
rect 233 164 253 166
rect 229 163 253 164
rect 3 156 257 157
rect 3 154 10 156
rect 12 154 50 156
rect 52 154 60 156
rect 62 154 91 156
rect 93 154 144 156
rect 146 154 155 156
rect 157 154 165 156
rect 167 154 196 156
rect 198 154 249 156
rect 251 154 257 156
rect 3 144 257 154
rect 3 142 10 144
rect 12 142 50 144
rect 52 142 60 144
rect 62 142 91 144
rect 93 142 144 144
rect 146 142 155 144
rect 157 142 165 144
rect 167 142 196 144
rect 198 142 249 144
rect 251 142 257 144
rect 3 141 257 142
rect 47 132 59 136
rect 47 130 49 132
rect 51 130 59 132
rect 124 134 148 135
rect 7 127 12 129
rect 7 125 9 127
rect 11 125 12 127
rect 7 123 12 125
rect 7 118 11 123
rect 7 116 8 118
rect 10 116 11 118
rect 7 104 11 116
rect 39 119 43 128
rect 47 119 51 130
rect 124 132 126 134
rect 128 132 148 134
rect 124 131 148 132
rect 7 102 9 104
rect 7 97 11 102
rect 7 95 9 97
rect 22 118 51 119
rect 22 116 26 118
rect 28 116 51 118
rect 22 115 51 116
rect 22 109 36 111
rect 38 109 43 111
rect 22 107 43 109
rect 39 101 43 107
rect 39 99 40 101
rect 42 99 43 101
rect 39 98 43 99
rect 47 110 51 115
rect 71 127 76 128
rect 71 125 72 127
rect 74 125 76 127
rect 71 119 76 125
rect 47 108 52 110
rect 47 106 49 108
rect 51 106 52 108
rect 47 101 52 106
rect 47 99 49 101
rect 51 99 52 101
rect 62 118 76 119
rect 62 116 66 118
rect 68 116 76 118
rect 62 115 76 116
rect 96 127 109 128
rect 96 125 99 127
rect 101 125 109 127
rect 96 123 109 125
rect 144 127 148 131
rect 96 122 106 123
rect 104 121 106 122
rect 108 121 109 123
rect 88 111 93 112
rect 70 110 83 111
rect 87 110 93 111
rect 70 108 76 110
rect 78 108 90 110
rect 92 108 93 110
rect 70 107 93 108
rect 79 105 93 107
rect 104 114 109 121
rect 144 125 145 127
rect 147 125 148 127
rect 47 97 52 99
rect 7 91 20 95
rect 7 90 11 91
rect 79 98 83 105
rect 88 96 93 105
rect 88 90 100 96
rect 144 103 148 125
rect 132 101 148 103
rect 132 99 134 101
rect 136 99 148 101
rect 132 98 148 99
rect 152 132 164 136
rect 152 130 154 132
rect 156 130 164 132
rect 229 134 253 135
rect 152 110 156 130
rect 229 132 231 134
rect 233 132 253 134
rect 229 131 253 132
rect 176 127 181 128
rect 176 125 177 127
rect 179 125 181 127
rect 176 119 181 125
rect 152 108 157 110
rect 152 106 154 108
rect 156 106 157 108
rect 152 101 157 106
rect 152 99 154 101
rect 156 99 157 101
rect 167 118 181 119
rect 167 116 171 118
rect 173 116 181 118
rect 167 115 181 116
rect 201 127 214 128
rect 201 125 204 127
rect 206 125 214 127
rect 201 123 214 125
rect 201 122 211 123
rect 209 121 211 122
rect 213 121 214 123
rect 193 111 198 112
rect 175 110 188 111
rect 192 110 198 111
rect 175 108 181 110
rect 183 108 195 110
rect 197 108 198 110
rect 175 107 198 108
rect 184 105 198 107
rect 209 114 214 121
rect 152 97 157 99
rect 184 101 188 105
rect 184 99 185 101
rect 187 99 188 101
rect 184 98 188 99
rect 193 96 198 105
rect 193 90 205 96
rect 249 103 253 131
rect 237 101 253 103
rect 237 99 239 101
rect 241 99 253 101
rect 237 98 253 99
rect 3 84 257 85
rect 3 82 10 84
rect 12 82 50 84
rect 52 82 124 84
rect 126 82 155 84
rect 157 82 229 84
rect 231 82 257 84
rect 3 72 257 82
rect 3 70 10 72
rect 12 70 50 72
rect 52 70 124 72
rect 126 70 155 72
rect 157 70 229 72
rect 231 70 257 72
rect 3 69 257 70
rect 7 63 11 64
rect 7 59 20 63
rect 7 57 9 59
rect 7 52 11 57
rect 7 50 9 52
rect 7 48 11 50
rect 39 55 43 56
rect 39 53 40 55
rect 42 53 43 55
rect 7 46 8 48
rect 10 46 11 48
rect 7 31 11 46
rect 39 47 43 53
rect 22 45 43 47
rect 22 43 36 45
rect 38 43 43 45
rect 47 55 52 57
rect 47 53 49 55
rect 51 53 52 55
rect 88 58 100 64
rect 47 48 52 53
rect 47 46 49 48
rect 51 46 52 48
rect 47 44 52 46
rect 47 39 51 44
rect 7 29 12 31
rect 7 27 9 29
rect 11 27 12 29
rect 7 25 12 27
rect 22 38 51 39
rect 22 36 26 38
rect 28 36 51 38
rect 22 35 51 36
rect 39 26 43 35
rect 47 24 51 35
rect 79 49 83 56
rect 88 49 93 58
rect 79 47 93 49
rect 70 46 93 47
rect 70 44 76 46
rect 78 44 90 46
rect 92 44 93 46
rect 70 43 83 44
rect 87 43 93 44
rect 88 42 93 43
rect 62 38 76 39
rect 62 36 66 38
rect 68 36 76 38
rect 62 35 76 36
rect 47 22 49 24
rect 51 22 59 24
rect 47 18 59 22
rect 71 29 76 35
rect 71 27 72 29
rect 74 27 76 29
rect 71 26 76 27
rect 104 33 109 40
rect 132 55 148 56
rect 132 53 134 55
rect 136 53 148 55
rect 132 51 148 53
rect 104 32 106 33
rect 96 31 106 32
rect 108 31 109 33
rect 96 29 109 31
rect 96 27 99 29
rect 101 27 109 29
rect 96 26 109 27
rect 144 29 148 51
rect 144 27 145 29
rect 147 27 148 29
rect 144 23 148 27
rect 124 22 148 23
rect 124 20 126 22
rect 128 20 148 22
rect 124 19 148 20
rect 152 55 157 57
rect 152 53 154 55
rect 156 53 157 55
rect 193 58 205 64
rect 152 48 157 53
rect 152 46 154 48
rect 156 46 157 48
rect 152 44 157 46
rect 152 24 156 44
rect 184 49 188 56
rect 193 49 198 58
rect 184 47 198 49
rect 175 46 198 47
rect 175 44 181 46
rect 183 44 195 46
rect 197 44 198 46
rect 175 43 188 44
rect 192 43 198 44
rect 193 42 198 43
rect 167 38 181 39
rect 167 36 171 38
rect 173 36 181 38
rect 167 35 181 36
rect 152 22 154 24
rect 156 22 164 24
rect 152 18 164 22
rect 176 29 181 35
rect 176 27 177 29
rect 179 27 181 29
rect 176 26 181 27
rect 209 33 214 40
rect 237 55 253 56
rect 237 53 239 55
rect 241 53 253 55
rect 237 51 253 53
rect 209 32 211 33
rect 201 31 211 32
rect 213 31 214 33
rect 201 29 214 31
rect 201 27 204 29
rect 206 27 214 29
rect 201 26 214 27
rect 249 23 253 51
rect 229 22 253 23
rect 229 20 231 22
rect 233 20 253 22
rect 229 19 253 20
rect 3 12 257 13
rect 3 10 10 12
rect 12 10 50 12
rect 52 10 60 12
rect 62 10 91 12
rect 93 10 144 12
rect 146 10 155 12
rect 157 10 165 12
rect 167 10 196 12
rect 198 10 249 12
rect 251 10 257 12
rect 3 5 257 10
<< alu2 >>
rect 71 271 104 272
rect 71 269 72 271
rect 74 269 99 271
rect 101 269 104 271
rect 71 268 104 269
rect 144 271 209 272
rect 144 269 145 271
rect 147 269 177 271
rect 179 269 204 271
rect 206 269 209 271
rect 144 268 209 269
rect 184 246 188 248
rect 39 245 157 246
rect 39 243 40 245
rect 42 243 154 245
rect 156 243 157 245
rect 39 242 157 243
rect 184 244 185 246
rect 187 244 188 246
rect 184 223 188 244
rect 7 219 188 223
rect 7 207 11 219
rect 7 205 8 207
rect 10 205 11 207
rect 7 198 11 205
rect 39 199 157 200
rect 39 197 40 199
rect 42 197 154 199
rect 156 197 157 199
rect 39 196 157 197
rect 130 190 184 191
rect 130 188 176 190
rect 178 188 184 190
rect 130 186 184 188
rect 71 173 104 174
rect 71 171 72 173
rect 74 171 99 173
rect 101 171 104 173
rect 71 170 104 171
rect 130 164 135 186
rect 144 173 209 174
rect 144 171 145 173
rect 147 171 177 173
rect 179 171 204 173
rect 206 171 209 173
rect 144 170 209 171
rect 7 160 135 164
rect 7 118 11 160
rect 71 127 104 128
rect 71 125 72 127
rect 74 125 99 127
rect 101 125 104 127
rect 71 124 104 125
rect 144 127 209 128
rect 144 125 145 127
rect 147 125 177 127
rect 179 125 204 127
rect 206 125 209 127
rect 144 124 209 125
rect 7 116 8 118
rect 10 116 11 118
rect 7 115 11 116
rect 39 101 157 102
rect 39 99 40 101
rect 42 99 154 101
rect 156 99 157 101
rect 39 98 157 99
rect 184 101 188 103
rect 184 99 185 101
rect 187 99 188 101
rect 184 78 188 99
rect 7 74 188 78
rect 7 48 11 74
rect 39 55 157 56
rect 39 53 40 55
rect 42 53 154 55
rect 156 53 157 55
rect 39 52 157 53
rect 7 46 8 48
rect 10 46 11 48
rect 7 45 11 46
rect 71 29 104 30
rect 71 27 72 29
rect 74 27 99 29
rect 101 27 104 29
rect 71 26 104 27
rect 144 29 209 30
rect 144 27 145 29
rect 147 27 177 29
rect 179 27 204 29
rect 206 27 209 29
rect 144 26 209 27
<< ptie >>
rect 8 288 14 290
rect 8 286 10 288
rect 12 286 14 288
rect 48 288 54 290
rect 48 286 50 288
rect 52 286 54 288
rect 8 284 14 286
rect 48 284 54 286
rect 89 288 95 290
rect 89 286 91 288
rect 93 286 95 288
rect 89 284 95 286
rect 153 288 159 290
rect 153 286 155 288
rect 157 286 159 288
rect 153 284 159 286
rect 194 288 200 290
rect 194 286 196 288
rect 198 286 200 288
rect 194 284 200 286
rect 8 156 14 158
rect 48 156 54 158
rect 8 154 10 156
rect 12 154 14 156
rect 8 152 14 154
rect 48 154 50 156
rect 52 154 54 156
rect 48 152 54 154
rect 89 156 95 158
rect 89 154 91 156
rect 93 154 95 156
rect 89 152 95 154
rect 153 156 159 158
rect 153 154 155 156
rect 157 154 159 156
rect 153 152 159 154
rect 194 156 200 158
rect 194 154 196 156
rect 198 154 200 156
rect 194 152 200 154
rect 8 144 14 146
rect 8 142 10 144
rect 12 142 14 144
rect 48 144 54 146
rect 48 142 50 144
rect 52 142 54 144
rect 8 140 14 142
rect 48 140 54 142
rect 89 144 95 146
rect 89 142 91 144
rect 93 142 95 144
rect 89 140 95 142
rect 153 144 159 146
rect 153 142 155 144
rect 157 142 159 144
rect 153 140 159 142
rect 194 144 200 146
rect 194 142 196 144
rect 198 142 200 144
rect 194 140 200 142
rect 8 12 14 14
rect 48 12 54 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 48 10 50 12
rect 52 10 54 12
rect 48 8 54 10
rect 89 12 95 14
rect 89 10 91 12
rect 93 10 95 12
rect 89 8 95 10
rect 153 12 159 14
rect 153 10 155 12
rect 157 10 159 12
rect 153 8 159 10
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
<< ntie >>
rect 8 228 14 230
rect 8 226 10 228
rect 12 226 14 228
rect 48 228 54 230
rect 8 224 14 226
rect 48 226 50 228
rect 52 226 54 228
rect 122 228 128 230
rect 48 224 54 226
rect 122 226 124 228
rect 126 226 128 228
rect 153 228 159 230
rect 122 224 128 226
rect 153 226 155 228
rect 157 226 159 228
rect 227 228 233 230
rect 153 224 159 226
rect 227 226 229 228
rect 231 226 233 228
rect 227 224 233 226
rect 8 216 14 218
rect 8 214 10 216
rect 12 214 14 216
rect 48 216 54 218
rect 8 212 14 214
rect 48 214 50 216
rect 52 214 54 216
rect 122 216 128 218
rect 48 212 54 214
rect 122 214 124 216
rect 126 214 128 216
rect 153 216 159 218
rect 122 212 128 214
rect 153 214 155 216
rect 157 214 159 216
rect 227 216 233 218
rect 153 212 159 214
rect 227 214 229 216
rect 231 214 233 216
rect 227 212 233 214
rect 8 84 14 86
rect 8 82 10 84
rect 12 82 14 84
rect 48 84 54 86
rect 8 80 14 82
rect 48 82 50 84
rect 52 82 54 84
rect 122 84 128 86
rect 48 80 54 82
rect 122 82 124 84
rect 126 82 128 84
rect 153 84 159 86
rect 122 80 128 82
rect 153 82 155 84
rect 157 82 159 84
rect 227 84 233 86
rect 153 80 159 82
rect 227 82 229 84
rect 231 82 233 84
rect 227 80 233 82
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 48 72 54 74
rect 8 68 14 70
rect 48 70 50 72
rect 52 70 54 72
rect 122 72 128 74
rect 48 68 54 70
rect 122 70 124 72
rect 126 70 128 72
rect 153 72 159 74
rect 122 68 128 70
rect 153 70 155 72
rect 157 70 159 72
rect 227 72 233 74
rect 153 68 159 70
rect 227 70 229 72
rect 231 70 233 72
rect 227 68 233 70
<< nmos >>
rect 14 267 16 276
rect 24 267 26 273
rect 34 267 36 273
rect 54 269 56 278
rect 67 269 69 280
rect 74 269 76 280
rect 95 267 97 276
rect 111 272 113 281
rect 121 272 123 281
rect 131 272 133 284
rect 138 272 140 284
rect 159 269 161 278
rect 172 269 174 280
rect 179 269 181 280
rect 200 267 202 276
rect 216 272 218 281
rect 226 272 228 281
rect 236 272 238 284
rect 243 272 245 284
rect 14 166 16 175
rect 24 169 26 175
rect 34 169 36 175
rect 54 164 56 173
rect 67 162 69 173
rect 74 162 76 173
rect 95 166 97 175
rect 111 161 113 170
rect 121 161 123 170
rect 131 158 133 170
rect 138 158 140 170
rect 159 164 161 173
rect 172 162 174 173
rect 179 162 181 173
rect 200 166 202 175
rect 216 161 218 170
rect 226 161 228 170
rect 236 158 238 170
rect 243 158 245 170
rect 14 123 16 132
rect 24 123 26 129
rect 34 123 36 129
rect 54 125 56 134
rect 67 125 69 136
rect 74 125 76 136
rect 95 123 97 132
rect 111 128 113 137
rect 121 128 123 137
rect 131 128 133 140
rect 138 128 140 140
rect 159 125 161 134
rect 172 125 174 136
rect 179 125 181 136
rect 200 123 202 132
rect 216 128 218 137
rect 226 128 228 137
rect 236 128 238 140
rect 243 128 245 140
rect 14 22 16 31
rect 24 25 26 31
rect 34 25 36 31
rect 54 20 56 29
rect 67 18 69 29
rect 74 18 76 29
rect 95 22 97 31
rect 111 17 113 26
rect 121 17 123 26
rect 131 14 133 26
rect 138 14 140 26
rect 159 20 161 29
rect 172 18 174 29
rect 179 18 181 29
rect 200 22 202 31
rect 216 17 218 26
rect 226 17 228 26
rect 236 14 238 26
rect 243 14 245 26
<< pmos >>
rect 14 237 16 255
rect 27 227 29 248
rect 34 227 36 248
rect 54 236 56 254
rect 64 234 66 247
rect 74 234 76 247
rect 103 227 105 254
rect 119 236 121 254
rect 129 236 131 254
rect 139 227 141 254
rect 159 236 161 254
rect 169 234 171 247
rect 179 234 181 247
rect 208 227 210 254
rect 224 236 226 254
rect 234 236 236 254
rect 244 227 246 254
rect 14 187 16 205
rect 27 194 29 215
rect 34 194 36 215
rect 54 188 56 206
rect 64 195 66 208
rect 74 195 76 208
rect 103 188 105 215
rect 119 188 121 206
rect 129 188 131 206
rect 139 188 141 215
rect 159 188 161 206
rect 169 195 171 208
rect 179 195 181 208
rect 208 188 210 215
rect 224 188 226 206
rect 234 188 236 206
rect 244 188 246 215
rect 14 93 16 111
rect 27 83 29 104
rect 34 83 36 104
rect 54 92 56 110
rect 64 90 66 103
rect 74 90 76 103
rect 103 83 105 110
rect 119 92 121 110
rect 129 92 131 110
rect 139 83 141 110
rect 159 92 161 110
rect 169 90 171 103
rect 179 90 181 103
rect 208 83 210 110
rect 224 92 226 110
rect 234 92 236 110
rect 244 83 246 110
rect 14 43 16 61
rect 27 50 29 71
rect 34 50 36 71
rect 54 44 56 62
rect 64 51 66 64
rect 74 51 76 64
rect 103 44 105 71
rect 119 44 121 62
rect 129 44 131 62
rect 139 44 141 71
rect 159 44 161 62
rect 169 51 171 64
rect 179 51 181 64
rect 208 44 210 71
rect 224 44 226 62
rect 234 44 236 62
rect 244 44 246 71
<< polyct0 >>
rect 16 260 18 262
rect 56 260 58 262
rect 127 260 129 262
rect 137 259 139 261
rect 161 260 163 262
rect 232 260 234 262
rect 242 259 244 261
rect 16 180 18 182
rect 56 180 58 182
rect 127 180 129 182
rect 137 181 139 183
rect 161 180 163 182
rect 232 180 234 182
rect 242 181 244 183
rect 16 116 18 118
rect 56 116 58 118
rect 127 116 129 118
rect 137 115 139 117
rect 161 116 163 118
rect 232 116 234 118
rect 242 115 244 117
rect 16 36 18 38
rect 56 36 58 38
rect 127 36 129 38
rect 137 37 139 39
rect 161 36 163 38
rect 232 36 234 38
rect 242 37 244 39
<< polyct1 >>
rect 26 260 28 262
rect 66 260 68 262
rect 36 253 38 255
rect 106 265 108 267
rect 76 252 78 254
rect 171 260 173 262
rect 90 252 92 254
rect 211 265 213 267
rect 181 252 183 254
rect 195 252 197 254
rect 36 187 38 189
rect 26 180 28 182
rect 76 188 78 190
rect 90 188 92 190
rect 66 180 68 182
rect 181 188 183 190
rect 195 188 197 190
rect 106 175 108 177
rect 171 180 173 182
rect 211 175 213 177
rect 26 116 28 118
rect 66 116 68 118
rect 36 109 38 111
rect 106 121 108 123
rect 76 108 78 110
rect 171 116 173 118
rect 90 108 92 110
rect 211 121 213 123
rect 181 108 183 110
rect 195 108 197 110
rect 36 43 38 45
rect 26 36 28 38
rect 76 44 78 46
rect 90 44 92 46
rect 66 36 68 38
rect 181 44 183 46
rect 195 44 197 46
rect 106 31 108 33
rect 171 36 173 38
rect 211 31 213 33
<< ndifct0 >>
rect 20 282 22 284
rect 39 282 41 284
rect 29 269 31 271
rect 79 276 81 278
rect 104 277 106 279
rect 90 269 92 271
rect 116 274 118 276
rect 184 276 186 278
rect 209 277 211 279
rect 195 269 197 271
rect 221 274 223 276
rect 29 171 31 173
rect 20 158 22 160
rect 90 171 92 173
rect 79 164 81 166
rect 104 163 106 165
rect 39 158 41 160
rect 116 166 118 168
rect 195 171 197 173
rect 184 164 186 166
rect 209 163 211 165
rect 221 166 223 168
rect 20 138 22 140
rect 39 138 41 140
rect 29 125 31 127
rect 79 132 81 134
rect 104 133 106 135
rect 90 125 92 127
rect 116 130 118 132
rect 184 132 186 134
rect 209 133 211 135
rect 195 125 197 127
rect 221 130 223 132
rect 29 27 31 29
rect 20 14 22 16
rect 90 27 92 29
rect 79 20 81 22
rect 104 19 106 21
rect 39 14 41 16
rect 116 22 118 24
rect 195 27 197 29
rect 184 20 186 22
rect 209 19 211 21
rect 221 22 223 24
<< ndifct1 >>
rect 60 286 62 288
rect 9 269 11 271
rect 144 286 146 288
rect 165 286 167 288
rect 49 274 51 276
rect 126 276 128 278
rect 249 286 251 288
rect 154 274 156 276
rect 231 276 233 278
rect 9 171 11 173
rect 49 166 51 168
rect 126 164 128 166
rect 60 154 62 156
rect 154 166 156 168
rect 144 154 146 156
rect 231 164 233 166
rect 165 154 167 156
rect 249 154 251 156
rect 60 142 62 144
rect 9 125 11 127
rect 144 142 146 144
rect 165 142 167 144
rect 49 130 51 132
rect 126 132 128 134
rect 249 142 251 144
rect 154 130 156 132
rect 231 132 233 134
rect 9 27 11 29
rect 49 22 51 24
rect 126 20 128 22
rect 60 10 62 12
rect 154 22 156 24
rect 144 10 146 12
rect 231 20 233 22
rect 165 10 167 12
rect 249 10 251 12
<< ntiect1 >>
rect 10 226 12 228
rect 50 226 52 228
rect 124 226 126 228
rect 155 226 157 228
rect 229 226 231 228
rect 10 214 12 216
rect 50 214 52 216
rect 124 214 126 216
rect 155 214 157 216
rect 229 214 231 216
rect 10 82 12 84
rect 50 82 52 84
rect 124 82 126 84
rect 155 82 157 84
rect 229 82 231 84
rect 10 70 12 72
rect 50 70 52 72
rect 124 70 126 72
rect 155 70 157 72
rect 229 70 231 72
<< ptiect1 >>
rect 10 286 12 288
rect 50 286 52 288
rect 91 286 93 288
rect 155 286 157 288
rect 196 286 198 288
rect 10 154 12 156
rect 50 154 52 156
rect 91 154 93 156
rect 155 154 157 156
rect 196 154 198 156
rect 10 142 12 144
rect 50 142 52 144
rect 91 142 93 144
rect 155 142 157 144
rect 196 142 198 144
rect 10 10 12 12
rect 50 10 52 12
rect 91 10 93 12
rect 155 10 157 12
rect 196 10 198 12
<< pdifct0 >>
rect 20 229 22 231
rect 39 236 41 238
rect 98 250 100 252
rect 59 238 61 240
rect 69 243 71 245
rect 69 236 71 238
rect 79 236 81 238
rect 108 236 110 238
rect 124 250 126 252
rect 124 243 126 245
rect 108 229 110 231
rect 144 235 146 237
rect 203 250 205 252
rect 164 238 166 240
rect 174 243 176 245
rect 174 236 176 238
rect 184 236 186 238
rect 213 236 215 238
rect 229 250 231 252
rect 229 243 231 245
rect 213 229 215 231
rect 249 235 251 237
rect 20 211 22 213
rect 39 204 41 206
rect 59 202 61 204
rect 69 204 71 206
rect 69 197 71 199
rect 79 204 81 206
rect 98 190 100 192
rect 108 211 110 213
rect 108 204 110 206
rect 124 197 126 199
rect 124 190 126 192
rect 144 205 146 207
rect 164 202 166 204
rect 174 204 176 206
rect 174 197 176 199
rect 184 204 186 206
rect 203 190 205 192
rect 213 211 215 213
rect 213 204 215 206
rect 229 197 231 199
rect 229 190 231 192
rect 249 205 251 207
rect 20 85 22 87
rect 39 92 41 94
rect 98 106 100 108
rect 59 94 61 96
rect 69 99 71 101
rect 69 92 71 94
rect 79 92 81 94
rect 108 92 110 94
rect 124 106 126 108
rect 124 99 126 101
rect 108 85 110 87
rect 144 91 146 93
rect 203 106 205 108
rect 164 94 166 96
rect 174 99 176 101
rect 174 92 176 94
rect 184 92 186 94
rect 213 92 215 94
rect 229 106 231 108
rect 229 99 231 101
rect 213 85 215 87
rect 249 91 251 93
rect 20 67 22 69
rect 39 60 41 62
rect 59 58 61 60
rect 69 60 71 62
rect 69 53 71 55
rect 79 60 81 62
rect 98 46 100 48
rect 108 67 110 69
rect 108 60 110 62
rect 124 53 126 55
rect 124 46 126 48
rect 144 61 146 63
rect 164 58 166 60
rect 174 60 176 62
rect 174 53 176 55
rect 184 60 186 62
rect 203 46 205 48
rect 213 67 215 69
rect 213 60 215 62
rect 229 53 231 55
rect 229 46 231 48
rect 249 61 251 63
<< pdifct1 >>
rect 9 246 11 248
rect 9 239 11 241
rect 49 250 51 252
rect 49 243 51 245
rect 134 243 136 245
rect 154 250 156 252
rect 154 243 156 245
rect 239 243 241 245
rect 9 201 11 203
rect 9 194 11 196
rect 49 197 51 199
rect 49 190 51 192
rect 134 197 136 199
rect 154 197 156 199
rect 154 190 156 192
rect 239 197 241 199
rect 9 102 11 104
rect 9 95 11 97
rect 49 106 51 108
rect 49 99 51 101
rect 134 99 136 101
rect 154 106 156 108
rect 154 99 156 101
rect 239 99 241 101
rect 9 57 11 59
rect 9 50 11 52
rect 49 53 51 55
rect 49 46 51 48
rect 134 53 136 55
rect 154 53 156 55
rect 154 46 156 48
rect 239 53 241 55
<< alu0 >>
rect 18 284 24 285
rect 18 282 20 284
rect 22 282 24 284
rect 18 281 24 282
rect 37 284 43 285
rect 37 282 39 284
rect 41 282 43 284
rect 37 281 43 282
rect 102 279 108 285
rect 63 278 83 279
rect 63 276 79 278
rect 81 276 83 278
rect 102 277 104 279
rect 106 277 108 279
rect 102 276 108 277
rect 115 276 119 278
rect 63 275 83 276
rect 15 271 33 272
rect 15 269 29 271
rect 31 269 33 271
rect 15 268 33 269
rect 15 262 19 268
rect 51 272 52 274
rect 63 271 67 275
rect 115 274 116 276
rect 118 274 119 276
rect 15 260 16 262
rect 18 260 19 262
rect 11 239 12 250
rect 15 247 19 260
rect 34 255 40 256
rect 15 243 30 247
rect 26 239 30 243
rect 55 267 67 271
rect 55 262 59 267
rect 55 260 56 262
rect 58 260 59 262
rect 55 248 59 260
rect 89 271 93 273
rect 89 269 90 271
rect 92 269 93 271
rect 89 263 93 269
rect 115 271 119 274
rect 115 267 139 271
rect 89 259 100 263
rect 96 253 100 259
rect 135 263 139 267
rect 115 262 131 263
rect 115 260 127 262
rect 129 260 131 262
rect 115 259 131 260
rect 135 261 140 263
rect 135 259 137 261
rect 139 259 140 261
rect 115 253 119 259
rect 135 257 140 259
rect 135 255 139 257
rect 96 252 119 253
rect 96 250 98 252
rect 100 250 119 252
rect 96 249 119 250
rect 55 245 72 248
rect 55 244 69 245
rect 68 243 69 244
rect 71 243 72 245
rect 57 240 63 241
rect 26 238 43 239
rect 26 236 39 238
rect 41 236 43 238
rect 26 235 43 236
rect 57 238 59 240
rect 61 238 63 240
rect 18 231 24 232
rect 18 229 20 231
rect 22 229 24 231
rect 57 229 63 238
rect 68 238 72 243
rect 68 236 69 238
rect 71 236 72 238
rect 68 234 72 236
rect 77 238 83 239
rect 77 236 79 238
rect 81 236 83 238
rect 77 229 83 236
rect 107 238 111 240
rect 107 236 108 238
rect 110 236 111 238
rect 107 231 111 236
rect 115 238 119 249
rect 123 252 139 255
rect 123 250 124 252
rect 126 251 139 252
rect 126 250 127 251
rect 123 245 127 250
rect 123 243 124 245
rect 126 243 127 245
rect 123 241 127 243
rect 207 279 213 285
rect 168 278 188 279
rect 168 276 184 278
rect 186 276 188 278
rect 207 277 209 279
rect 211 277 213 279
rect 207 276 213 277
rect 220 276 224 278
rect 168 275 188 276
rect 156 272 157 274
rect 168 271 172 275
rect 220 274 221 276
rect 223 274 224 276
rect 160 267 172 271
rect 160 262 164 267
rect 160 260 161 262
rect 163 260 164 262
rect 160 248 164 260
rect 194 271 198 273
rect 194 269 195 271
rect 197 269 198 271
rect 194 263 198 269
rect 220 271 224 274
rect 220 267 244 271
rect 194 259 205 263
rect 201 253 205 259
rect 240 263 244 267
rect 220 262 236 263
rect 220 260 232 262
rect 234 260 236 262
rect 220 259 236 260
rect 240 261 245 263
rect 240 259 242 261
rect 244 259 245 261
rect 220 253 224 259
rect 240 257 245 259
rect 240 255 244 257
rect 201 252 224 253
rect 201 250 203 252
rect 205 250 224 252
rect 201 249 224 250
rect 160 245 177 248
rect 160 244 174 245
rect 173 243 174 244
rect 176 243 177 245
rect 162 240 168 241
rect 162 238 164 240
rect 166 238 168 240
rect 115 237 148 238
rect 115 235 144 237
rect 146 235 148 237
rect 115 234 148 235
rect 107 229 108 231
rect 110 229 111 231
rect 162 229 168 238
rect 173 238 177 243
rect 173 236 174 238
rect 176 236 177 238
rect 173 234 177 236
rect 182 238 188 239
rect 182 236 184 238
rect 186 236 188 238
rect 182 229 188 236
rect 212 238 216 240
rect 212 236 213 238
rect 215 236 216 238
rect 212 231 216 236
rect 220 238 224 249
rect 228 252 244 255
rect 228 250 229 252
rect 231 251 244 252
rect 231 250 232 251
rect 228 245 232 250
rect 228 243 229 245
rect 231 243 232 245
rect 228 241 232 243
rect 220 237 253 238
rect 220 235 249 237
rect 251 235 253 237
rect 220 234 253 235
rect 212 229 213 231
rect 215 229 216 231
rect 18 211 20 213
rect 22 211 24 213
rect 18 210 24 211
rect 26 206 43 207
rect 26 204 39 206
rect 41 204 43 206
rect 26 203 43 204
rect 57 204 63 213
rect 11 192 12 203
rect 26 199 30 203
rect 57 202 59 204
rect 61 202 63 204
rect 57 201 63 202
rect 68 206 72 208
rect 68 204 69 206
rect 71 204 72 206
rect 15 195 30 199
rect 15 182 19 195
rect 68 199 72 204
rect 77 206 83 213
rect 107 211 108 213
rect 110 211 111 213
rect 77 204 79 206
rect 81 204 83 206
rect 77 203 83 204
rect 107 206 111 211
rect 107 204 108 206
rect 110 204 111 206
rect 107 202 111 204
rect 115 207 148 208
rect 115 205 144 207
rect 146 205 148 207
rect 115 204 148 205
rect 162 204 168 213
rect 68 198 69 199
rect 55 197 69 198
rect 71 197 72 199
rect 55 194 72 197
rect 34 186 40 187
rect 15 180 16 182
rect 18 180 19 182
rect 15 174 19 180
rect 15 173 33 174
rect 15 171 29 173
rect 31 171 33 173
rect 15 170 33 171
rect 55 182 59 194
rect 115 193 119 204
rect 162 202 164 204
rect 166 202 168 204
rect 162 201 168 202
rect 173 206 177 208
rect 173 204 174 206
rect 176 204 177 206
rect 96 192 119 193
rect 96 190 98 192
rect 100 190 119 192
rect 96 189 119 190
rect 96 183 100 189
rect 55 180 56 182
rect 58 180 59 182
rect 55 175 59 180
rect 55 171 67 175
rect 51 168 52 170
rect 63 167 67 171
rect 89 179 100 183
rect 89 173 93 179
rect 115 183 119 189
rect 123 199 127 201
rect 123 197 124 199
rect 126 197 127 199
rect 123 192 127 197
rect 123 190 124 192
rect 126 191 127 192
rect 126 190 139 191
rect 123 187 139 190
rect 135 185 139 187
rect 135 183 140 185
rect 115 182 131 183
rect 115 180 127 182
rect 129 180 131 182
rect 115 179 131 180
rect 135 181 137 183
rect 139 181 140 183
rect 135 179 140 181
rect 89 171 90 173
rect 92 171 93 173
rect 89 169 93 171
rect 135 175 139 179
rect 115 171 139 175
rect 115 168 119 171
rect 63 166 83 167
rect 115 166 116 168
rect 118 166 119 168
rect 63 164 79 166
rect 81 164 83 166
rect 63 163 83 164
rect 102 165 108 166
rect 102 163 104 165
rect 106 163 108 165
rect 115 164 119 166
rect 173 199 177 204
rect 182 206 188 213
rect 212 211 213 213
rect 215 211 216 213
rect 182 204 184 206
rect 186 204 188 206
rect 182 203 188 204
rect 212 206 216 211
rect 212 204 213 206
rect 215 204 216 206
rect 212 202 216 204
rect 220 207 253 208
rect 220 205 249 207
rect 251 205 253 207
rect 220 204 253 205
rect 173 198 174 199
rect 160 197 174 198
rect 176 197 177 199
rect 160 194 177 197
rect 160 182 164 194
rect 220 193 224 204
rect 201 192 224 193
rect 201 190 203 192
rect 205 190 224 192
rect 201 189 224 190
rect 201 183 205 189
rect 160 180 161 182
rect 163 180 164 182
rect 160 175 164 180
rect 160 171 172 175
rect 156 168 157 170
rect 18 160 24 161
rect 18 158 20 160
rect 22 158 24 160
rect 18 157 24 158
rect 37 160 43 161
rect 37 158 39 160
rect 41 158 43 160
rect 37 157 43 158
rect 102 157 108 163
rect 168 167 172 171
rect 194 179 205 183
rect 194 173 198 179
rect 220 183 224 189
rect 228 199 232 201
rect 228 197 229 199
rect 231 197 232 199
rect 228 192 232 197
rect 228 190 229 192
rect 231 191 232 192
rect 231 190 244 191
rect 228 187 244 190
rect 240 185 244 187
rect 240 183 245 185
rect 220 182 236 183
rect 220 180 232 182
rect 234 180 236 182
rect 220 179 236 180
rect 240 181 242 183
rect 244 181 245 183
rect 240 179 245 181
rect 194 171 195 173
rect 197 171 198 173
rect 194 169 198 171
rect 240 175 244 179
rect 220 171 244 175
rect 220 168 224 171
rect 168 166 188 167
rect 220 166 221 168
rect 223 166 224 168
rect 168 164 184 166
rect 186 164 188 166
rect 168 163 188 164
rect 207 165 213 166
rect 207 163 209 165
rect 211 163 213 165
rect 220 164 224 166
rect 207 157 213 163
rect 18 140 24 141
rect 18 138 20 140
rect 22 138 24 140
rect 18 137 24 138
rect 37 140 43 141
rect 37 138 39 140
rect 41 138 43 140
rect 37 137 43 138
rect 102 135 108 141
rect 63 134 83 135
rect 63 132 79 134
rect 81 132 83 134
rect 102 133 104 135
rect 106 133 108 135
rect 102 132 108 133
rect 115 132 119 134
rect 63 131 83 132
rect 15 127 33 128
rect 15 125 29 127
rect 31 125 33 127
rect 15 124 33 125
rect 15 118 19 124
rect 51 128 52 130
rect 63 127 67 131
rect 115 130 116 132
rect 118 130 119 132
rect 15 116 16 118
rect 18 116 19 118
rect 11 95 12 106
rect 15 103 19 116
rect 34 111 40 112
rect 15 99 30 103
rect 26 95 30 99
rect 55 123 67 127
rect 55 118 59 123
rect 55 116 56 118
rect 58 116 59 118
rect 55 104 59 116
rect 89 127 93 129
rect 89 125 90 127
rect 92 125 93 127
rect 89 119 93 125
rect 115 127 119 130
rect 115 123 139 127
rect 89 115 100 119
rect 96 109 100 115
rect 135 119 139 123
rect 115 118 131 119
rect 115 116 127 118
rect 129 116 131 118
rect 115 115 131 116
rect 135 117 140 119
rect 135 115 137 117
rect 139 115 140 117
rect 115 109 119 115
rect 135 113 140 115
rect 135 111 139 113
rect 96 108 119 109
rect 96 106 98 108
rect 100 106 119 108
rect 96 105 119 106
rect 55 101 72 104
rect 55 100 69 101
rect 68 99 69 100
rect 71 99 72 101
rect 57 96 63 97
rect 26 94 43 95
rect 26 92 39 94
rect 41 92 43 94
rect 26 91 43 92
rect 57 94 59 96
rect 61 94 63 96
rect 18 87 24 88
rect 18 85 20 87
rect 22 85 24 87
rect 57 85 63 94
rect 68 94 72 99
rect 68 92 69 94
rect 71 92 72 94
rect 68 90 72 92
rect 77 94 83 95
rect 77 92 79 94
rect 81 92 83 94
rect 77 85 83 92
rect 107 94 111 96
rect 107 92 108 94
rect 110 92 111 94
rect 107 87 111 92
rect 115 94 119 105
rect 123 108 139 111
rect 123 106 124 108
rect 126 107 139 108
rect 126 106 127 107
rect 123 101 127 106
rect 123 99 124 101
rect 126 99 127 101
rect 123 97 127 99
rect 207 135 213 141
rect 168 134 188 135
rect 168 132 184 134
rect 186 132 188 134
rect 207 133 209 135
rect 211 133 213 135
rect 207 132 213 133
rect 220 132 224 134
rect 168 131 188 132
rect 156 128 157 130
rect 168 127 172 131
rect 220 130 221 132
rect 223 130 224 132
rect 160 123 172 127
rect 160 118 164 123
rect 160 116 161 118
rect 163 116 164 118
rect 160 104 164 116
rect 194 127 198 129
rect 194 125 195 127
rect 197 125 198 127
rect 194 119 198 125
rect 220 127 224 130
rect 220 123 244 127
rect 194 115 205 119
rect 201 109 205 115
rect 240 119 244 123
rect 220 118 236 119
rect 220 116 232 118
rect 234 116 236 118
rect 220 115 236 116
rect 240 117 245 119
rect 240 115 242 117
rect 244 115 245 117
rect 220 109 224 115
rect 240 113 245 115
rect 240 111 244 113
rect 201 108 224 109
rect 201 106 203 108
rect 205 106 224 108
rect 201 105 224 106
rect 160 101 177 104
rect 160 100 174 101
rect 173 99 174 100
rect 176 99 177 101
rect 162 96 168 97
rect 162 94 164 96
rect 166 94 168 96
rect 115 93 148 94
rect 115 91 144 93
rect 146 91 148 93
rect 115 90 148 91
rect 107 85 108 87
rect 110 85 111 87
rect 162 85 168 94
rect 173 94 177 99
rect 173 92 174 94
rect 176 92 177 94
rect 173 90 177 92
rect 182 94 188 95
rect 182 92 184 94
rect 186 92 188 94
rect 182 85 188 92
rect 212 94 216 96
rect 212 92 213 94
rect 215 92 216 94
rect 212 87 216 92
rect 220 94 224 105
rect 228 108 244 111
rect 228 106 229 108
rect 231 107 244 108
rect 231 106 232 107
rect 228 101 232 106
rect 228 99 229 101
rect 231 99 232 101
rect 228 97 232 99
rect 220 93 253 94
rect 220 91 249 93
rect 251 91 253 93
rect 220 90 253 91
rect 212 85 213 87
rect 215 85 216 87
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 26 62 43 63
rect 26 60 39 62
rect 41 60 43 62
rect 26 59 43 60
rect 57 60 63 69
rect 11 48 12 59
rect 26 55 30 59
rect 57 58 59 60
rect 61 58 63 60
rect 57 57 63 58
rect 68 62 72 64
rect 68 60 69 62
rect 71 60 72 62
rect 15 51 30 55
rect 15 38 19 51
rect 68 55 72 60
rect 77 62 83 69
rect 107 67 108 69
rect 110 67 111 69
rect 77 60 79 62
rect 81 60 83 62
rect 77 59 83 60
rect 107 62 111 67
rect 107 60 108 62
rect 110 60 111 62
rect 107 58 111 60
rect 115 63 148 64
rect 115 61 144 63
rect 146 61 148 63
rect 115 60 148 61
rect 162 60 168 69
rect 68 54 69 55
rect 55 53 69 54
rect 71 53 72 55
rect 55 50 72 53
rect 34 42 40 43
rect 15 36 16 38
rect 18 36 19 38
rect 15 30 19 36
rect 15 29 33 30
rect 15 27 29 29
rect 31 27 33 29
rect 15 26 33 27
rect 55 38 59 50
rect 115 49 119 60
rect 162 58 164 60
rect 166 58 168 60
rect 162 57 168 58
rect 173 62 177 64
rect 173 60 174 62
rect 176 60 177 62
rect 96 48 119 49
rect 96 46 98 48
rect 100 46 119 48
rect 96 45 119 46
rect 96 39 100 45
rect 55 36 56 38
rect 58 36 59 38
rect 55 31 59 36
rect 55 27 67 31
rect 51 24 52 26
rect 63 23 67 27
rect 89 35 100 39
rect 89 29 93 35
rect 115 39 119 45
rect 123 55 127 57
rect 123 53 124 55
rect 126 53 127 55
rect 123 48 127 53
rect 123 46 124 48
rect 126 47 127 48
rect 126 46 139 47
rect 123 43 139 46
rect 135 41 139 43
rect 135 39 140 41
rect 115 38 131 39
rect 115 36 127 38
rect 129 36 131 38
rect 115 35 131 36
rect 135 37 137 39
rect 139 37 140 39
rect 135 35 140 37
rect 89 27 90 29
rect 92 27 93 29
rect 89 25 93 27
rect 135 31 139 35
rect 115 27 139 31
rect 115 24 119 27
rect 63 22 83 23
rect 115 22 116 24
rect 118 22 119 24
rect 63 20 79 22
rect 81 20 83 22
rect 63 19 83 20
rect 102 21 108 22
rect 102 19 104 21
rect 106 19 108 21
rect 115 20 119 22
rect 173 55 177 60
rect 182 62 188 69
rect 212 67 213 69
rect 215 67 216 69
rect 182 60 184 62
rect 186 60 188 62
rect 182 59 188 60
rect 212 62 216 67
rect 212 60 213 62
rect 215 60 216 62
rect 212 58 216 60
rect 220 63 253 64
rect 220 61 249 63
rect 251 61 253 63
rect 220 60 253 61
rect 173 54 174 55
rect 160 53 174 54
rect 176 53 177 55
rect 160 50 177 53
rect 160 38 164 50
rect 220 49 224 60
rect 201 48 224 49
rect 201 46 203 48
rect 205 46 224 48
rect 201 45 224 46
rect 201 39 205 45
rect 160 36 161 38
rect 163 36 164 38
rect 160 31 164 36
rect 160 27 172 31
rect 156 24 157 26
rect 18 16 24 17
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 37 16 43 17
rect 37 14 39 16
rect 41 14 43 16
rect 37 13 43 14
rect 102 13 108 19
rect 168 23 172 27
rect 194 35 205 39
rect 194 29 198 35
rect 220 39 224 45
rect 228 55 232 57
rect 228 53 229 55
rect 231 53 232 55
rect 228 48 232 53
rect 228 46 229 48
rect 231 47 232 48
rect 231 46 244 47
rect 228 43 244 46
rect 240 41 244 43
rect 240 39 245 41
rect 220 38 236 39
rect 220 36 232 38
rect 234 36 236 38
rect 220 35 236 36
rect 240 37 242 39
rect 244 37 245 39
rect 240 35 245 37
rect 194 27 195 29
rect 197 27 198 29
rect 194 25 198 27
rect 240 31 244 35
rect 220 27 244 31
rect 220 24 224 27
rect 168 22 188 23
rect 220 22 221 24
rect 223 22 224 24
rect 168 20 184 22
rect 186 20 188 22
rect 168 19 188 20
rect 207 21 213 22
rect 207 19 209 21
rect 211 19 213 21
rect 220 20 224 22
rect 207 13 213 19
<< via1 >>
rect 40 243 42 245
rect 72 269 74 271
rect 99 269 101 271
rect 145 269 147 271
rect 177 269 179 271
rect 154 243 156 245
rect 204 269 206 271
rect 185 244 187 246
rect 8 205 10 207
rect 40 197 42 199
rect 72 171 74 173
rect 99 171 101 173
rect 145 171 147 173
rect 154 197 156 199
rect 176 188 178 190
rect 177 171 179 173
rect 204 171 206 173
rect 8 116 10 118
rect 40 99 42 101
rect 72 125 74 127
rect 99 125 101 127
rect 145 125 147 127
rect 177 125 179 127
rect 154 99 156 101
rect 204 125 206 127
rect 185 99 187 101
rect 40 53 42 55
rect 8 46 10 48
rect 72 27 74 29
rect 99 27 101 29
rect 145 27 147 29
rect 154 53 156 55
rect 177 27 179 29
rect 204 27 206 29
<< labels >>
rlabel alu1 89 73 89 73 1 Vdd
rlabel alu1 65 73 65 73 6 vdd
rlabel alu1 87 8 87 8 1 Vss
rlabel alu1 194 73 194 73 1 Vdd
rlabel alu1 170 73 170 73 6 vdd
rlabel alu1 192 8 192 8 1 Vss
rlabel alu1 186 53 186 53 1 cin
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 89 81 89 81 5 Vdd
rlabel alu1 65 81 65 81 8 vdd
rlabel alu1 87 146 87 146 5 Vss
rlabel alu1 194 81 194 81 5 Vdd
rlabel alu1 170 81 170 81 8 vdd
rlabel alu1 192 146 192 146 5 Vss
rlabel alu1 25 81 25 81 8 vdd
rlabel alu1 25 217 25 217 6 vdd
rlabel alu1 192 152 192 152 1 Vss
rlabel alu1 170 217 170 217 6 vdd
rlabel alu1 194 217 194 217 1 Vdd
rlabel alu1 87 152 87 152 1 Vss
rlabel alu1 65 217 65 217 6 vdd
rlabel alu1 89 217 89 217 1 Vdd
rlabel alu1 9 254 9 254 5 cout
rlabel alu1 25 225 25 225 8 vdd
rlabel alu1 192 290 192 290 5 Vss
rlabel alu1 170 225 170 225 8 vdd
rlabel alu1 194 225 194 225 5 Vdd
rlabel alu1 87 290 87 290 5 Vss
rlabel alu1 65 225 65 225 8 vdd
rlabel alu1 89 225 89 225 5 Vdd
rlabel alu1 9 110 9 110 1 cout1
rlabel alu1 9 44 9 44 1 cout0
rlabel alu1 9 188 9 188 1 cout2
rlabel alu1 98 61 98 61 1 b0
rlabel alu1 73 33 73 33 1 a0
rlabel alu1 107 36 107 36 1 a0
rlabel alu1 98 93 98 93 1 b1
rlabel alu1 107 118 107 118 1 a1
rlabel alu1 73 121 73 121 1 a1
rlabel alu1 98 205 98 205 1 b2
rlabel alu1 73 177 73 177 1 a2
rlabel alu1 107 180 107 180 1 a2
rlabel alu1 98 237 98 237 1 b3
rlabel alu1 73 265 73 265 1 a3
rlabel alu1 107 262 107 262 1 a3
rlabel alu1 251 40 251 40 1 s0
rlabel alu1 251 114 251 114 1 s1
rlabel alu1 251 184 251 184 1 s2
rlabel alu1 251 258 251 258 1 s3
<< end >>
