magic
tech scmos
timestamp 1607850035
<< ab >>
rect 88 293 94 298
rect 202 293 208 298
rect 4 5 44 293
rect 53 261 157 293
rect 53 229 93 261
rect 94 229 157 261
rect 46 213 51 229
rect 53 213 157 229
rect 53 181 93 213
rect 94 181 157 213
rect 53 117 157 181
rect 53 85 93 117
rect 94 85 157 117
rect 46 69 51 85
rect 53 69 157 85
rect 53 37 93 69
rect 94 37 157 69
rect 53 5 157 37
rect 167 261 271 293
rect 272 285 276 293
rect 167 229 207 261
rect 208 229 271 261
rect 167 213 271 229
rect 272 213 274 229
rect 167 181 207 213
rect 208 181 271 213
rect 167 117 271 181
rect 272 141 276 157
rect 167 85 207 117
rect 208 85 271 117
rect 167 69 271 85
rect 272 69 274 85
rect 167 37 207 69
rect 208 37 271 69
rect 167 5 271 37
rect 272 5 276 13
rect 278 5 318 293
rect 319 285 383 293
rect 322 229 383 285
rect 319 213 383 229
rect 322 157 383 213
rect 319 141 383 157
rect 322 85 383 141
rect 319 69 383 85
rect 322 13 383 69
rect 319 5 383 13
rect 387 5 451 293
rect 455 5 518 293
rect 520 285 560 293
rect 562 285 632 293
rect 521 229 560 285
rect 563 229 626 285
rect 520 213 560 229
rect 561 213 626 229
rect 627 213 632 229
rect 521 157 560 213
rect 563 157 626 213
rect 520 141 560 157
rect 562 141 632 157
rect 521 85 560 141
rect 563 85 626 141
rect 520 69 560 85
rect 561 69 626 85
rect 627 69 632 85
rect 521 13 560 69
rect 563 13 626 69
rect 520 5 560 13
rect 562 5 632 13
rect 88 0 94 5
rect 202 0 208 5
<< nwell >>
rect -1 181 632 261
rect -1 37 632 117
<< pwell >>
rect -1 261 632 298
rect -1 117 632 181
rect -1 0 632 37
<< poly >>
rect 13 276 15 281
rect 23 273 25 278
rect 33 273 35 278
rect 62 278 64 282
rect 75 280 77 285
rect 82 280 84 285
rect 105 289 130 291
rect 105 281 107 289
rect 118 281 120 285
rect 128 281 130 289
rect 138 284 140 289
rect 145 284 147 289
rect 102 279 107 281
rect 102 276 104 279
rect 13 264 15 267
rect 23 264 25 267
rect 13 262 19 264
rect 13 260 15 262
rect 17 260 19 262
rect 13 258 19 260
rect 23 262 29 264
rect 23 260 25 262
rect 27 260 29 262
rect 23 258 29 260
rect 13 255 15 258
rect 26 248 28 258
rect 33 257 35 267
rect 62 264 64 269
rect 75 264 77 269
rect 62 262 68 264
rect 62 260 64 262
rect 66 260 68 262
rect 62 258 68 260
rect 72 262 78 264
rect 72 260 74 262
rect 76 260 78 262
rect 72 258 78 260
rect 33 255 39 257
rect 33 253 35 255
rect 37 253 39 255
rect 62 254 64 258
rect 33 251 39 253
rect 33 248 35 251
rect 13 232 15 237
rect 72 247 74 258
rect 82 256 84 269
rect 176 278 178 282
rect 189 280 191 285
rect 196 280 198 285
rect 219 289 244 291
rect 219 281 221 289
rect 232 281 234 285
rect 242 281 244 289
rect 252 284 254 289
rect 259 284 261 289
rect 118 269 120 272
rect 111 267 120 269
rect 128 268 130 272
rect 138 269 140 272
rect 102 259 104 267
rect 111 265 113 267
rect 115 265 120 267
rect 111 263 120 265
rect 136 267 140 269
rect 136 264 138 267
rect 118 259 120 263
rect 132 262 138 264
rect 145 263 147 272
rect 216 279 221 281
rect 216 276 218 279
rect 176 264 178 269
rect 189 264 191 269
rect 132 260 134 262
rect 136 260 138 262
rect 99 257 112 259
rect 118 257 128 259
rect 132 258 138 260
rect 99 256 101 257
rect 82 254 88 256
rect 82 252 84 254
rect 86 252 88 254
rect 82 250 88 252
rect 95 254 101 256
rect 110 254 112 257
rect 126 254 128 257
rect 136 254 138 258
rect 142 261 148 263
rect 142 259 144 261
rect 146 259 148 261
rect 142 257 148 259
rect 146 254 148 257
rect 176 262 182 264
rect 176 260 178 262
rect 180 260 182 262
rect 176 258 182 260
rect 186 262 192 264
rect 186 260 188 262
rect 190 260 192 262
rect 186 258 192 260
rect 176 254 178 258
rect 95 252 97 254
rect 99 252 101 254
rect 95 250 101 252
rect 82 247 84 250
rect 62 232 64 236
rect 72 229 74 234
rect 82 229 84 234
rect 26 223 28 227
rect 33 223 35 227
rect 126 232 128 236
rect 136 232 138 236
rect 110 223 112 227
rect 186 247 188 258
rect 196 256 198 269
rect 287 280 289 285
rect 294 280 296 285
rect 329 289 348 291
rect 232 269 234 272
rect 225 267 234 269
rect 242 268 244 272
rect 252 269 254 272
rect 216 259 218 267
rect 225 265 227 267
rect 229 265 234 267
rect 225 263 234 265
rect 250 267 254 269
rect 250 264 252 267
rect 232 259 234 263
rect 246 262 252 264
rect 259 263 261 272
rect 307 278 309 282
rect 329 279 331 289
rect 339 281 341 285
rect 346 281 348 289
rect 423 289 442 291
rect 356 281 358 286
rect 363 281 365 286
rect 373 281 375 286
rect 396 281 398 286
rect 406 281 408 286
rect 413 281 415 286
rect 423 281 425 289
rect 430 281 432 285
rect 246 260 248 262
rect 250 260 252 262
rect 213 257 226 259
rect 232 257 242 259
rect 246 258 252 260
rect 213 256 215 257
rect 196 254 202 256
rect 196 252 198 254
rect 200 252 202 254
rect 196 250 202 252
rect 209 254 215 256
rect 224 254 226 257
rect 240 254 242 257
rect 250 254 252 258
rect 256 261 262 263
rect 256 259 258 261
rect 260 259 262 261
rect 256 257 262 259
rect 260 254 262 257
rect 287 256 289 269
rect 294 264 296 269
rect 307 264 309 269
rect 293 262 299 264
rect 293 260 295 262
rect 297 260 299 262
rect 293 258 299 260
rect 303 262 309 264
rect 303 260 305 262
rect 307 260 309 262
rect 303 258 309 260
rect 283 254 289 256
rect 209 252 211 254
rect 213 252 215 254
rect 209 250 215 252
rect 196 247 198 250
rect 176 232 178 236
rect 186 229 188 234
rect 196 229 198 234
rect 146 223 148 227
rect 240 232 242 236
rect 250 232 252 236
rect 224 223 226 227
rect 283 252 285 254
rect 287 252 289 254
rect 283 250 289 252
rect 287 247 289 250
rect 297 247 299 258
rect 307 254 309 258
rect 329 255 331 273
rect 339 264 341 273
rect 335 262 341 264
rect 335 260 337 262
rect 339 260 341 262
rect 335 258 341 260
rect 346 260 348 273
rect 356 270 358 273
rect 352 268 358 270
rect 352 266 354 268
rect 356 266 358 268
rect 352 264 358 266
rect 346 258 358 260
rect 363 259 365 273
rect 440 279 442 289
rect 490 289 509 291
rect 463 281 465 286
rect 473 281 475 286
rect 480 281 482 286
rect 490 281 492 289
rect 497 281 499 285
rect 373 269 375 272
rect 396 269 398 272
rect 370 267 376 269
rect 370 265 372 267
rect 374 265 376 267
rect 370 263 376 265
rect 395 267 401 269
rect 395 265 397 267
rect 399 265 401 267
rect 395 263 401 265
rect 329 244 331 247
rect 322 242 331 244
rect 339 243 341 258
rect 345 252 351 254
rect 345 250 347 252
rect 349 250 351 252
rect 345 248 351 250
rect 346 243 348 248
rect 356 243 358 258
rect 362 257 368 259
rect 362 255 364 257
rect 366 255 368 257
rect 362 253 368 255
rect 363 243 365 253
rect 373 245 375 263
rect 396 245 398 263
rect 406 259 408 273
rect 413 270 415 273
rect 413 268 419 270
rect 413 266 415 268
rect 417 266 419 268
rect 413 264 419 266
rect 423 260 425 273
rect 403 257 409 259
rect 403 255 405 257
rect 407 255 409 257
rect 403 253 409 255
rect 413 258 425 260
rect 430 264 432 273
rect 430 262 436 264
rect 430 260 432 262
rect 434 260 436 262
rect 430 258 436 260
rect 322 240 324 242
rect 326 240 328 242
rect 322 238 328 240
rect 287 229 289 234
rect 297 229 299 234
rect 307 232 309 236
rect 260 223 262 227
rect 406 243 408 253
rect 413 243 415 258
rect 420 252 426 254
rect 420 250 422 252
rect 424 250 426 252
rect 420 248 426 250
rect 423 243 425 248
rect 430 243 432 258
rect 440 255 442 273
rect 507 279 509 289
rect 589 289 614 291
rect 529 276 531 281
rect 463 269 465 272
rect 462 267 468 269
rect 462 265 464 267
rect 466 265 468 267
rect 462 263 468 265
rect 440 244 442 247
rect 463 245 465 263
rect 473 259 475 273
rect 480 270 482 273
rect 480 268 486 270
rect 480 266 482 268
rect 484 266 486 268
rect 480 264 486 266
rect 490 260 492 273
rect 470 257 476 259
rect 470 255 472 257
rect 474 255 476 257
rect 470 253 476 255
rect 480 258 492 260
rect 497 264 499 273
rect 497 262 503 264
rect 497 260 499 262
rect 501 260 503 262
rect 497 258 503 260
rect 440 242 449 244
rect 443 240 445 242
rect 447 240 449 242
rect 443 238 449 240
rect 473 243 475 253
rect 480 243 482 258
rect 487 252 493 254
rect 487 250 489 252
rect 491 250 493 252
rect 487 248 493 250
rect 490 243 492 248
rect 497 243 499 258
rect 507 255 509 273
rect 539 273 541 278
rect 549 273 551 278
rect 572 284 574 289
rect 579 284 581 289
rect 589 281 591 289
rect 599 281 601 285
rect 612 281 614 289
rect 612 279 617 281
rect 615 276 617 279
rect 529 264 531 267
rect 539 264 541 267
rect 529 262 535 264
rect 529 260 531 262
rect 533 260 535 262
rect 529 258 535 260
rect 539 262 545 264
rect 539 260 541 262
rect 543 260 545 262
rect 539 258 545 260
rect 529 255 531 258
rect 507 244 509 247
rect 507 242 516 244
rect 510 240 512 242
rect 514 240 516 242
rect 510 238 516 240
rect 542 248 544 258
rect 549 257 551 267
rect 572 263 574 272
rect 579 269 581 272
rect 579 267 583 269
rect 589 268 591 272
rect 599 269 601 272
rect 581 264 583 267
rect 599 267 608 269
rect 599 265 604 267
rect 606 265 608 267
rect 571 261 577 263
rect 571 259 573 261
rect 575 259 577 261
rect 571 257 577 259
rect 581 262 587 264
rect 581 260 583 262
rect 585 260 587 262
rect 581 258 587 260
rect 599 263 608 265
rect 599 259 601 263
rect 615 259 617 267
rect 549 255 555 257
rect 549 253 551 255
rect 553 253 555 255
rect 571 254 573 257
rect 581 254 583 258
rect 591 257 601 259
rect 607 257 620 259
rect 591 254 593 257
rect 607 254 609 257
rect 618 256 620 257
rect 618 254 624 256
rect 549 251 555 253
rect 549 248 551 251
rect 529 232 531 237
rect 339 223 341 227
rect 346 223 348 227
rect 356 223 358 227
rect 363 223 365 227
rect 373 223 375 227
rect 396 223 398 227
rect 406 223 408 227
rect 413 223 415 227
rect 423 223 425 227
rect 430 223 432 227
rect 463 223 465 227
rect 473 223 475 227
rect 480 223 482 227
rect 490 223 492 227
rect 497 223 499 227
rect 581 232 583 236
rect 591 232 593 236
rect 542 223 544 227
rect 549 223 551 227
rect 571 223 573 227
rect 618 252 620 254
rect 622 252 624 254
rect 618 250 624 252
rect 607 223 609 227
rect 26 215 28 219
rect 33 215 35 219
rect 13 205 15 210
rect 110 215 112 219
rect 62 206 64 210
rect 72 208 74 213
rect 82 208 84 213
rect 13 184 15 187
rect 26 184 28 194
rect 33 191 35 194
rect 33 189 39 191
rect 33 187 35 189
rect 37 187 39 189
rect 33 185 39 187
rect 13 182 19 184
rect 13 180 15 182
rect 17 180 19 182
rect 13 178 19 180
rect 23 182 29 184
rect 23 180 25 182
rect 27 180 29 182
rect 23 178 29 180
rect 13 175 15 178
rect 23 175 25 178
rect 33 175 35 185
rect 62 184 64 188
rect 72 184 74 195
rect 82 192 84 195
rect 82 190 88 192
rect 82 188 84 190
rect 86 188 88 190
rect 82 186 88 188
rect 95 190 101 192
rect 95 188 97 190
rect 99 188 101 190
rect 146 215 148 219
rect 126 206 128 210
rect 136 206 138 210
rect 224 215 226 219
rect 176 206 178 210
rect 186 208 188 213
rect 196 208 198 213
rect 95 186 101 188
rect 62 182 68 184
rect 62 180 64 182
rect 66 180 68 182
rect 62 178 68 180
rect 72 182 78 184
rect 72 180 74 182
rect 76 180 78 182
rect 72 178 78 180
rect 62 173 64 178
rect 75 173 77 178
rect 82 173 84 186
rect 99 185 101 186
rect 110 185 112 188
rect 126 185 128 188
rect 99 183 112 185
rect 118 183 128 185
rect 136 184 138 188
rect 146 185 148 188
rect 102 175 104 183
rect 118 179 120 183
rect 111 177 120 179
rect 132 182 138 184
rect 132 180 134 182
rect 136 180 138 182
rect 132 178 138 180
rect 142 183 148 185
rect 142 181 144 183
rect 146 181 148 183
rect 142 179 148 181
rect 176 184 178 188
rect 186 184 188 195
rect 196 192 198 195
rect 196 190 202 192
rect 196 188 198 190
rect 200 188 202 190
rect 196 186 202 188
rect 209 190 215 192
rect 209 188 211 190
rect 213 188 215 190
rect 260 215 262 219
rect 240 206 242 210
rect 250 206 252 210
rect 339 215 341 219
rect 346 215 348 219
rect 356 215 358 219
rect 363 215 365 219
rect 373 215 375 219
rect 396 215 398 219
rect 406 215 408 219
rect 413 215 415 219
rect 423 215 425 219
rect 430 215 432 219
rect 463 215 465 219
rect 473 215 475 219
rect 480 215 482 219
rect 490 215 492 219
rect 497 215 499 219
rect 287 208 289 213
rect 297 208 299 213
rect 307 206 309 210
rect 287 192 289 195
rect 283 190 289 192
rect 283 188 285 190
rect 287 188 289 190
rect 209 186 215 188
rect 176 182 182 184
rect 176 180 178 182
rect 180 180 182 182
rect 111 175 113 177
rect 115 175 120 177
rect 13 161 15 166
rect 23 164 25 169
rect 33 164 35 169
rect 62 160 64 164
rect 111 173 120 175
rect 136 175 138 178
rect 118 170 120 173
rect 128 170 130 174
rect 136 173 140 175
rect 138 170 140 173
rect 145 170 147 179
rect 176 178 182 180
rect 186 182 192 184
rect 186 180 188 182
rect 190 180 192 182
rect 186 178 192 180
rect 176 173 178 178
rect 189 173 191 178
rect 196 173 198 186
rect 213 185 215 186
rect 224 185 226 188
rect 240 185 242 188
rect 213 183 226 185
rect 232 183 242 185
rect 250 184 252 188
rect 260 185 262 188
rect 283 186 289 188
rect 216 175 218 183
rect 232 179 234 183
rect 225 177 234 179
rect 246 182 252 184
rect 246 180 248 182
rect 250 180 252 182
rect 246 178 252 180
rect 256 183 262 185
rect 256 181 258 183
rect 260 181 262 183
rect 256 179 262 181
rect 225 175 227 177
rect 229 175 234 177
rect 102 163 104 166
rect 75 157 77 162
rect 82 157 84 162
rect 102 161 107 163
rect 105 153 107 161
rect 118 157 120 161
rect 128 153 130 161
rect 176 160 178 164
rect 225 173 234 175
rect 250 175 252 178
rect 232 170 234 173
rect 242 170 244 174
rect 250 173 254 175
rect 252 170 254 173
rect 259 170 261 179
rect 287 173 289 186
rect 297 184 299 195
rect 322 202 328 204
rect 322 200 324 202
rect 326 200 328 202
rect 322 198 331 200
rect 329 195 331 198
rect 307 184 309 188
rect 293 182 299 184
rect 293 180 295 182
rect 297 180 299 182
rect 293 178 299 180
rect 303 182 309 184
rect 303 180 305 182
rect 307 180 309 182
rect 303 178 309 180
rect 294 173 296 178
rect 307 173 309 178
rect 216 163 218 166
rect 138 153 140 158
rect 145 153 147 158
rect 105 151 130 153
rect 189 157 191 162
rect 196 157 198 162
rect 216 161 221 163
rect 219 153 221 161
rect 232 157 234 161
rect 242 153 244 161
rect 329 169 331 187
rect 339 184 341 199
rect 346 194 348 199
rect 345 192 351 194
rect 345 190 347 192
rect 349 190 351 192
rect 345 188 351 190
rect 356 184 358 199
rect 363 189 365 199
rect 443 202 449 204
rect 443 200 445 202
rect 447 200 449 202
rect 335 182 341 184
rect 335 180 337 182
rect 339 180 341 182
rect 335 178 341 180
rect 339 169 341 178
rect 346 182 358 184
rect 362 187 368 189
rect 362 185 364 187
rect 366 185 368 187
rect 362 183 368 185
rect 346 169 348 182
rect 352 176 358 178
rect 352 174 354 176
rect 356 174 358 176
rect 352 172 358 174
rect 356 169 358 172
rect 363 169 365 183
rect 373 179 375 197
rect 396 179 398 197
rect 406 189 408 199
rect 403 187 409 189
rect 403 185 405 187
rect 407 185 409 187
rect 403 183 409 185
rect 413 184 415 199
rect 423 194 425 199
rect 420 192 426 194
rect 420 190 422 192
rect 424 190 426 192
rect 420 188 426 190
rect 430 184 432 199
rect 440 198 449 200
rect 440 195 442 198
rect 542 215 544 219
rect 549 215 551 219
rect 571 215 573 219
rect 529 205 531 210
rect 510 202 516 204
rect 510 200 512 202
rect 514 200 516 202
rect 370 177 376 179
rect 370 175 372 177
rect 374 175 376 177
rect 370 173 376 175
rect 395 177 401 179
rect 395 175 397 177
rect 399 175 401 177
rect 395 173 401 175
rect 373 170 375 173
rect 396 170 398 173
rect 252 153 254 158
rect 259 153 261 158
rect 287 157 289 162
rect 294 157 296 162
rect 219 151 244 153
rect 307 160 309 164
rect 329 153 331 163
rect 406 169 408 183
rect 413 182 425 184
rect 413 176 419 178
rect 413 174 415 176
rect 417 174 419 176
rect 413 172 419 174
rect 413 169 415 172
rect 423 169 425 182
rect 430 182 436 184
rect 430 180 432 182
rect 434 180 436 182
rect 430 178 436 180
rect 430 169 432 178
rect 440 169 442 187
rect 463 179 465 197
rect 473 189 475 199
rect 470 187 476 189
rect 470 185 472 187
rect 474 185 476 187
rect 470 183 476 185
rect 480 184 482 199
rect 490 194 492 199
rect 487 192 493 194
rect 487 190 489 192
rect 491 190 493 192
rect 487 188 493 190
rect 497 184 499 199
rect 507 198 516 200
rect 507 195 509 198
rect 462 177 468 179
rect 462 175 464 177
rect 466 175 468 177
rect 462 173 468 175
rect 463 170 465 173
rect 339 157 341 161
rect 346 153 348 161
rect 356 156 358 161
rect 363 156 365 161
rect 373 156 375 161
rect 396 156 398 161
rect 406 156 408 161
rect 413 156 415 161
rect 329 151 348 153
rect 423 153 425 161
rect 430 157 432 161
rect 440 153 442 163
rect 473 169 475 183
rect 480 182 492 184
rect 480 176 486 178
rect 480 174 482 176
rect 484 174 486 176
rect 480 172 486 174
rect 480 169 482 172
rect 490 169 492 182
rect 497 182 503 184
rect 497 180 499 182
rect 501 180 503 182
rect 497 178 503 180
rect 497 169 499 178
rect 507 169 509 187
rect 529 184 531 187
rect 542 184 544 194
rect 549 191 551 194
rect 549 189 555 191
rect 549 187 551 189
rect 553 187 555 189
rect 607 215 609 219
rect 581 206 583 210
rect 591 206 593 210
rect 618 190 624 192
rect 618 188 620 190
rect 622 188 624 190
rect 549 185 555 187
rect 571 185 573 188
rect 529 182 535 184
rect 529 180 531 182
rect 533 180 535 182
rect 529 178 535 180
rect 539 182 545 184
rect 539 180 541 182
rect 543 180 545 182
rect 539 178 545 180
rect 529 175 531 178
rect 539 175 541 178
rect 549 175 551 185
rect 571 183 577 185
rect 571 181 573 183
rect 575 181 577 183
rect 571 179 577 181
rect 581 184 583 188
rect 591 185 593 188
rect 607 185 609 188
rect 618 186 624 188
rect 618 185 620 186
rect 581 182 587 184
rect 591 183 601 185
rect 607 183 620 185
rect 581 180 583 182
rect 585 180 587 182
rect 572 170 574 179
rect 581 178 587 180
rect 599 179 601 183
rect 581 175 583 178
rect 579 173 583 175
rect 599 177 608 179
rect 599 175 604 177
rect 606 175 608 177
rect 615 175 617 183
rect 579 170 581 173
rect 589 170 591 174
rect 599 173 608 175
rect 599 170 601 173
rect 463 156 465 161
rect 473 156 475 161
rect 480 156 482 161
rect 423 151 442 153
rect 490 153 492 161
rect 497 157 499 161
rect 507 153 509 163
rect 529 161 531 166
rect 539 164 541 169
rect 549 164 551 169
rect 490 151 509 153
rect 615 163 617 166
rect 612 161 617 163
rect 572 153 574 158
rect 579 153 581 158
rect 589 153 591 161
rect 599 157 601 161
rect 612 153 614 161
rect 589 151 614 153
rect 13 132 15 137
rect 23 129 25 134
rect 33 129 35 134
rect 62 134 64 138
rect 75 136 77 141
rect 82 136 84 141
rect 105 145 130 147
rect 105 137 107 145
rect 118 137 120 141
rect 128 137 130 145
rect 138 140 140 145
rect 145 140 147 145
rect 102 135 107 137
rect 102 132 104 135
rect 13 120 15 123
rect 23 120 25 123
rect 13 118 19 120
rect 13 116 15 118
rect 17 116 19 118
rect 13 114 19 116
rect 23 118 29 120
rect 23 116 25 118
rect 27 116 29 118
rect 23 114 29 116
rect 13 111 15 114
rect 26 104 28 114
rect 33 113 35 123
rect 62 120 64 125
rect 75 120 77 125
rect 62 118 68 120
rect 62 116 64 118
rect 66 116 68 118
rect 62 114 68 116
rect 72 118 78 120
rect 72 116 74 118
rect 76 116 78 118
rect 72 114 78 116
rect 33 111 39 113
rect 33 109 35 111
rect 37 109 39 111
rect 62 110 64 114
rect 33 107 39 109
rect 33 104 35 107
rect 13 88 15 93
rect 72 103 74 114
rect 82 112 84 125
rect 176 134 178 138
rect 189 136 191 141
rect 196 136 198 141
rect 219 145 244 147
rect 219 137 221 145
rect 232 137 234 141
rect 242 137 244 145
rect 252 140 254 145
rect 259 140 261 145
rect 118 125 120 128
rect 111 123 120 125
rect 128 124 130 128
rect 138 125 140 128
rect 102 115 104 123
rect 111 121 113 123
rect 115 121 120 123
rect 111 119 120 121
rect 136 123 140 125
rect 136 120 138 123
rect 118 115 120 119
rect 132 118 138 120
rect 145 119 147 128
rect 216 135 221 137
rect 216 132 218 135
rect 176 120 178 125
rect 189 120 191 125
rect 132 116 134 118
rect 136 116 138 118
rect 99 113 112 115
rect 118 113 128 115
rect 132 114 138 116
rect 99 112 101 113
rect 82 110 88 112
rect 82 108 84 110
rect 86 108 88 110
rect 82 106 88 108
rect 95 110 101 112
rect 110 110 112 113
rect 126 110 128 113
rect 136 110 138 114
rect 142 117 148 119
rect 142 115 144 117
rect 146 115 148 117
rect 142 113 148 115
rect 146 110 148 113
rect 176 118 182 120
rect 176 116 178 118
rect 180 116 182 118
rect 176 114 182 116
rect 186 118 192 120
rect 186 116 188 118
rect 190 116 192 118
rect 186 114 192 116
rect 176 110 178 114
rect 95 108 97 110
rect 99 108 101 110
rect 95 106 101 108
rect 82 103 84 106
rect 62 88 64 92
rect 72 85 74 90
rect 82 85 84 90
rect 26 79 28 83
rect 33 79 35 83
rect 126 88 128 92
rect 136 88 138 92
rect 110 79 112 83
rect 186 103 188 114
rect 196 112 198 125
rect 287 136 289 141
rect 294 136 296 141
rect 329 145 348 147
rect 232 125 234 128
rect 225 123 234 125
rect 242 124 244 128
rect 252 125 254 128
rect 216 115 218 123
rect 225 121 227 123
rect 229 121 234 123
rect 225 119 234 121
rect 250 123 254 125
rect 250 120 252 123
rect 232 115 234 119
rect 246 118 252 120
rect 259 119 261 128
rect 307 134 309 138
rect 329 135 331 145
rect 339 137 341 141
rect 346 137 348 145
rect 423 145 442 147
rect 356 137 358 142
rect 363 137 365 142
rect 373 137 375 142
rect 396 137 398 142
rect 406 137 408 142
rect 413 137 415 142
rect 423 137 425 145
rect 430 137 432 141
rect 246 116 248 118
rect 250 116 252 118
rect 213 113 226 115
rect 232 113 242 115
rect 246 114 252 116
rect 213 112 215 113
rect 196 110 202 112
rect 196 108 198 110
rect 200 108 202 110
rect 196 106 202 108
rect 209 110 215 112
rect 224 110 226 113
rect 240 110 242 113
rect 250 110 252 114
rect 256 117 262 119
rect 256 115 258 117
rect 260 115 262 117
rect 256 113 262 115
rect 260 110 262 113
rect 287 112 289 125
rect 294 120 296 125
rect 307 120 309 125
rect 293 118 299 120
rect 293 116 295 118
rect 297 116 299 118
rect 293 114 299 116
rect 303 118 309 120
rect 303 116 305 118
rect 307 116 309 118
rect 303 114 309 116
rect 283 110 289 112
rect 209 108 211 110
rect 213 108 215 110
rect 209 106 215 108
rect 196 103 198 106
rect 176 88 178 92
rect 186 85 188 90
rect 196 85 198 90
rect 146 79 148 83
rect 240 88 242 92
rect 250 88 252 92
rect 224 79 226 83
rect 283 108 285 110
rect 287 108 289 110
rect 283 106 289 108
rect 287 103 289 106
rect 297 103 299 114
rect 307 110 309 114
rect 329 111 331 129
rect 339 120 341 129
rect 335 118 341 120
rect 335 116 337 118
rect 339 116 341 118
rect 335 114 341 116
rect 346 116 348 129
rect 356 126 358 129
rect 352 124 358 126
rect 352 122 354 124
rect 356 122 358 124
rect 352 120 358 122
rect 346 114 358 116
rect 363 115 365 129
rect 440 135 442 145
rect 490 145 509 147
rect 463 137 465 142
rect 473 137 475 142
rect 480 137 482 142
rect 490 137 492 145
rect 497 137 499 141
rect 373 125 375 128
rect 396 125 398 128
rect 370 123 376 125
rect 370 121 372 123
rect 374 121 376 123
rect 370 119 376 121
rect 395 123 401 125
rect 395 121 397 123
rect 399 121 401 123
rect 395 119 401 121
rect 329 100 331 103
rect 322 98 331 100
rect 339 99 341 114
rect 345 108 351 110
rect 345 106 347 108
rect 349 106 351 108
rect 345 104 351 106
rect 346 99 348 104
rect 356 99 358 114
rect 362 113 368 115
rect 362 111 364 113
rect 366 111 368 113
rect 362 109 368 111
rect 363 99 365 109
rect 373 101 375 119
rect 396 101 398 119
rect 406 115 408 129
rect 413 126 415 129
rect 413 124 419 126
rect 413 122 415 124
rect 417 122 419 124
rect 413 120 419 122
rect 423 116 425 129
rect 403 113 409 115
rect 403 111 405 113
rect 407 111 409 113
rect 403 109 409 111
rect 413 114 425 116
rect 430 120 432 129
rect 430 118 436 120
rect 430 116 432 118
rect 434 116 436 118
rect 430 114 436 116
rect 322 96 324 98
rect 326 96 328 98
rect 322 94 328 96
rect 287 85 289 90
rect 297 85 299 90
rect 307 88 309 92
rect 260 79 262 83
rect 406 99 408 109
rect 413 99 415 114
rect 420 108 426 110
rect 420 106 422 108
rect 424 106 426 108
rect 420 104 426 106
rect 423 99 425 104
rect 430 99 432 114
rect 440 111 442 129
rect 507 135 509 145
rect 589 145 614 147
rect 529 132 531 137
rect 463 125 465 128
rect 462 123 468 125
rect 462 121 464 123
rect 466 121 468 123
rect 462 119 468 121
rect 440 100 442 103
rect 463 101 465 119
rect 473 115 475 129
rect 480 126 482 129
rect 480 124 486 126
rect 480 122 482 124
rect 484 122 486 124
rect 480 120 486 122
rect 490 116 492 129
rect 470 113 476 115
rect 470 111 472 113
rect 474 111 476 113
rect 470 109 476 111
rect 480 114 492 116
rect 497 120 499 129
rect 497 118 503 120
rect 497 116 499 118
rect 501 116 503 118
rect 497 114 503 116
rect 440 98 449 100
rect 443 96 445 98
rect 447 96 449 98
rect 443 94 449 96
rect 473 99 475 109
rect 480 99 482 114
rect 487 108 493 110
rect 487 106 489 108
rect 491 106 493 108
rect 487 104 493 106
rect 490 99 492 104
rect 497 99 499 114
rect 507 111 509 129
rect 539 129 541 134
rect 549 129 551 134
rect 572 140 574 145
rect 579 140 581 145
rect 589 137 591 145
rect 599 137 601 141
rect 612 137 614 145
rect 612 135 617 137
rect 615 132 617 135
rect 529 120 531 123
rect 539 120 541 123
rect 529 118 535 120
rect 529 116 531 118
rect 533 116 535 118
rect 529 114 535 116
rect 539 118 545 120
rect 539 116 541 118
rect 543 116 545 118
rect 539 114 545 116
rect 529 111 531 114
rect 507 100 509 103
rect 507 98 516 100
rect 510 96 512 98
rect 514 96 516 98
rect 510 94 516 96
rect 542 104 544 114
rect 549 113 551 123
rect 572 119 574 128
rect 579 125 581 128
rect 579 123 583 125
rect 589 124 591 128
rect 599 125 601 128
rect 581 120 583 123
rect 599 123 608 125
rect 599 121 604 123
rect 606 121 608 123
rect 571 117 577 119
rect 571 115 573 117
rect 575 115 577 117
rect 571 113 577 115
rect 581 118 587 120
rect 581 116 583 118
rect 585 116 587 118
rect 581 114 587 116
rect 599 119 608 121
rect 599 115 601 119
rect 615 115 617 123
rect 549 111 555 113
rect 549 109 551 111
rect 553 109 555 111
rect 571 110 573 113
rect 581 110 583 114
rect 591 113 601 115
rect 607 113 620 115
rect 591 110 593 113
rect 607 110 609 113
rect 618 112 620 113
rect 618 110 624 112
rect 549 107 555 109
rect 549 104 551 107
rect 529 88 531 93
rect 339 79 341 83
rect 346 79 348 83
rect 356 79 358 83
rect 363 79 365 83
rect 373 79 375 83
rect 396 79 398 83
rect 406 79 408 83
rect 413 79 415 83
rect 423 79 425 83
rect 430 79 432 83
rect 463 79 465 83
rect 473 79 475 83
rect 480 79 482 83
rect 490 79 492 83
rect 497 79 499 83
rect 581 88 583 92
rect 591 88 593 92
rect 542 79 544 83
rect 549 79 551 83
rect 571 79 573 83
rect 618 108 620 110
rect 622 108 624 110
rect 618 106 624 108
rect 607 79 609 83
rect 26 71 28 75
rect 33 71 35 75
rect 13 61 15 66
rect 110 71 112 75
rect 62 62 64 66
rect 72 64 74 69
rect 82 64 84 69
rect 13 40 15 43
rect 26 40 28 50
rect 33 47 35 50
rect 33 45 39 47
rect 33 43 35 45
rect 37 43 39 45
rect 33 41 39 43
rect 13 38 19 40
rect 13 36 15 38
rect 17 36 19 38
rect 13 34 19 36
rect 23 38 29 40
rect 23 36 25 38
rect 27 36 29 38
rect 23 34 29 36
rect 13 31 15 34
rect 23 31 25 34
rect 33 31 35 41
rect 62 40 64 44
rect 72 40 74 51
rect 82 48 84 51
rect 82 46 88 48
rect 82 44 84 46
rect 86 44 88 46
rect 82 42 88 44
rect 95 46 101 48
rect 95 44 97 46
rect 99 44 101 46
rect 146 71 148 75
rect 126 62 128 66
rect 136 62 138 66
rect 224 71 226 75
rect 176 62 178 66
rect 186 64 188 69
rect 196 64 198 69
rect 95 42 101 44
rect 62 38 68 40
rect 62 36 64 38
rect 66 36 68 38
rect 62 34 68 36
rect 72 38 78 40
rect 72 36 74 38
rect 76 36 78 38
rect 72 34 78 36
rect 62 29 64 34
rect 75 29 77 34
rect 82 29 84 42
rect 99 41 101 42
rect 110 41 112 44
rect 126 41 128 44
rect 99 39 112 41
rect 118 39 128 41
rect 136 40 138 44
rect 146 41 148 44
rect 102 31 104 39
rect 118 35 120 39
rect 111 33 120 35
rect 132 38 138 40
rect 132 36 134 38
rect 136 36 138 38
rect 132 34 138 36
rect 142 39 148 41
rect 142 37 144 39
rect 146 37 148 39
rect 142 35 148 37
rect 176 40 178 44
rect 186 40 188 51
rect 196 48 198 51
rect 196 46 202 48
rect 196 44 198 46
rect 200 44 202 46
rect 196 42 202 44
rect 209 46 215 48
rect 209 44 211 46
rect 213 44 215 46
rect 260 71 262 75
rect 240 62 242 66
rect 250 62 252 66
rect 339 71 341 75
rect 346 71 348 75
rect 356 71 358 75
rect 363 71 365 75
rect 373 71 375 75
rect 396 71 398 75
rect 406 71 408 75
rect 413 71 415 75
rect 423 71 425 75
rect 430 71 432 75
rect 463 71 465 75
rect 473 71 475 75
rect 480 71 482 75
rect 490 71 492 75
rect 497 71 499 75
rect 287 64 289 69
rect 297 64 299 69
rect 307 62 309 66
rect 287 48 289 51
rect 283 46 289 48
rect 283 44 285 46
rect 287 44 289 46
rect 209 42 215 44
rect 176 38 182 40
rect 176 36 178 38
rect 180 36 182 38
rect 111 31 113 33
rect 115 31 120 33
rect 13 17 15 22
rect 23 20 25 25
rect 33 20 35 25
rect 62 16 64 20
rect 111 29 120 31
rect 136 31 138 34
rect 118 26 120 29
rect 128 26 130 30
rect 136 29 140 31
rect 138 26 140 29
rect 145 26 147 35
rect 176 34 182 36
rect 186 38 192 40
rect 186 36 188 38
rect 190 36 192 38
rect 186 34 192 36
rect 176 29 178 34
rect 189 29 191 34
rect 196 29 198 42
rect 213 41 215 42
rect 224 41 226 44
rect 240 41 242 44
rect 213 39 226 41
rect 232 39 242 41
rect 250 40 252 44
rect 260 41 262 44
rect 283 42 289 44
rect 216 31 218 39
rect 232 35 234 39
rect 225 33 234 35
rect 246 38 252 40
rect 246 36 248 38
rect 250 36 252 38
rect 246 34 252 36
rect 256 39 262 41
rect 256 37 258 39
rect 260 37 262 39
rect 256 35 262 37
rect 225 31 227 33
rect 229 31 234 33
rect 102 19 104 22
rect 75 13 77 18
rect 82 13 84 18
rect 102 17 107 19
rect 105 9 107 17
rect 118 13 120 17
rect 128 9 130 17
rect 176 16 178 20
rect 225 29 234 31
rect 250 31 252 34
rect 232 26 234 29
rect 242 26 244 30
rect 250 29 254 31
rect 252 26 254 29
rect 259 26 261 35
rect 287 29 289 42
rect 297 40 299 51
rect 322 58 328 60
rect 322 56 324 58
rect 326 56 328 58
rect 322 54 331 56
rect 329 51 331 54
rect 307 40 309 44
rect 293 38 299 40
rect 293 36 295 38
rect 297 36 299 38
rect 293 34 299 36
rect 303 38 309 40
rect 303 36 305 38
rect 307 36 309 38
rect 303 34 309 36
rect 294 29 296 34
rect 307 29 309 34
rect 216 19 218 22
rect 138 9 140 14
rect 145 9 147 14
rect 105 7 130 9
rect 189 13 191 18
rect 196 13 198 18
rect 216 17 221 19
rect 219 9 221 17
rect 232 13 234 17
rect 242 9 244 17
rect 329 25 331 43
rect 339 40 341 55
rect 346 50 348 55
rect 345 48 351 50
rect 345 46 347 48
rect 349 46 351 48
rect 345 44 351 46
rect 356 40 358 55
rect 363 45 365 55
rect 443 58 449 60
rect 443 56 445 58
rect 447 56 449 58
rect 335 38 341 40
rect 335 36 337 38
rect 339 36 341 38
rect 335 34 341 36
rect 339 25 341 34
rect 346 38 358 40
rect 362 43 368 45
rect 362 41 364 43
rect 366 41 368 43
rect 362 39 368 41
rect 346 25 348 38
rect 352 32 358 34
rect 352 30 354 32
rect 356 30 358 32
rect 352 28 358 30
rect 356 25 358 28
rect 363 25 365 39
rect 373 35 375 53
rect 396 35 398 53
rect 406 45 408 55
rect 403 43 409 45
rect 403 41 405 43
rect 407 41 409 43
rect 403 39 409 41
rect 413 40 415 55
rect 423 50 425 55
rect 420 48 426 50
rect 420 46 422 48
rect 424 46 426 48
rect 420 44 426 46
rect 430 40 432 55
rect 440 54 449 56
rect 440 51 442 54
rect 542 71 544 75
rect 549 71 551 75
rect 571 71 573 75
rect 529 61 531 66
rect 510 58 516 60
rect 510 56 512 58
rect 514 56 516 58
rect 370 33 376 35
rect 370 31 372 33
rect 374 31 376 33
rect 370 29 376 31
rect 395 33 401 35
rect 395 31 397 33
rect 399 31 401 33
rect 395 29 401 31
rect 373 26 375 29
rect 396 26 398 29
rect 252 9 254 14
rect 259 9 261 14
rect 287 13 289 18
rect 294 13 296 18
rect 219 7 244 9
rect 307 16 309 20
rect 329 9 331 19
rect 406 25 408 39
rect 413 38 425 40
rect 413 32 419 34
rect 413 30 415 32
rect 417 30 419 32
rect 413 28 419 30
rect 413 25 415 28
rect 423 25 425 38
rect 430 38 436 40
rect 430 36 432 38
rect 434 36 436 38
rect 430 34 436 36
rect 430 25 432 34
rect 440 25 442 43
rect 463 35 465 53
rect 473 45 475 55
rect 470 43 476 45
rect 470 41 472 43
rect 474 41 476 43
rect 470 39 476 41
rect 480 40 482 55
rect 490 50 492 55
rect 487 48 493 50
rect 487 46 489 48
rect 491 46 493 48
rect 487 44 493 46
rect 497 40 499 55
rect 507 54 516 56
rect 507 51 509 54
rect 462 33 468 35
rect 462 31 464 33
rect 466 31 468 33
rect 462 29 468 31
rect 463 26 465 29
rect 339 13 341 17
rect 346 9 348 17
rect 356 12 358 17
rect 363 12 365 17
rect 373 12 375 17
rect 396 12 398 17
rect 406 12 408 17
rect 413 12 415 17
rect 329 7 348 9
rect 423 9 425 17
rect 430 13 432 17
rect 440 9 442 19
rect 473 25 475 39
rect 480 38 492 40
rect 480 32 486 34
rect 480 30 482 32
rect 484 30 486 32
rect 480 28 486 30
rect 480 25 482 28
rect 490 25 492 38
rect 497 38 503 40
rect 497 36 499 38
rect 501 36 503 38
rect 497 34 503 36
rect 497 25 499 34
rect 507 25 509 43
rect 529 40 531 43
rect 542 40 544 50
rect 549 47 551 50
rect 549 45 555 47
rect 549 43 551 45
rect 553 43 555 45
rect 607 71 609 75
rect 581 62 583 66
rect 591 62 593 66
rect 618 46 624 48
rect 618 44 620 46
rect 622 44 624 46
rect 549 41 555 43
rect 571 41 573 44
rect 529 38 535 40
rect 529 36 531 38
rect 533 36 535 38
rect 529 34 535 36
rect 539 38 545 40
rect 539 36 541 38
rect 543 36 545 38
rect 539 34 545 36
rect 529 31 531 34
rect 539 31 541 34
rect 549 31 551 41
rect 571 39 577 41
rect 571 37 573 39
rect 575 37 577 39
rect 571 35 577 37
rect 581 40 583 44
rect 591 41 593 44
rect 607 41 609 44
rect 618 42 624 44
rect 618 41 620 42
rect 581 38 587 40
rect 591 39 601 41
rect 607 39 620 41
rect 581 36 583 38
rect 585 36 587 38
rect 572 26 574 35
rect 581 34 587 36
rect 599 35 601 39
rect 581 31 583 34
rect 579 29 583 31
rect 599 33 608 35
rect 599 31 604 33
rect 606 31 608 33
rect 615 31 617 39
rect 579 26 581 29
rect 589 26 591 30
rect 599 29 608 31
rect 599 26 601 29
rect 463 12 465 17
rect 473 12 475 17
rect 480 12 482 17
rect 423 7 442 9
rect 490 9 492 17
rect 497 13 499 17
rect 507 9 509 19
rect 529 17 531 22
rect 539 20 541 25
rect 549 20 551 25
rect 490 7 509 9
rect 615 19 617 22
rect 612 17 617 19
rect 572 9 574 14
rect 579 9 581 14
rect 589 9 591 17
rect 599 13 601 17
rect 612 9 614 17
rect 589 7 614 9
<< ndif >>
rect 17 284 23 286
rect 17 282 19 284
rect 21 282 23 284
rect 17 280 23 282
rect 36 284 42 286
rect 66 288 73 290
rect 66 286 68 288
rect 70 286 73 288
rect 36 282 38 284
rect 40 282 42 284
rect 36 280 42 282
rect 17 276 21 280
rect 8 273 13 276
rect 6 271 13 273
rect 6 269 8 271
rect 10 269 13 271
rect 6 267 13 269
rect 15 273 21 276
rect 37 273 42 280
rect 66 280 73 286
rect 149 288 155 290
rect 149 286 151 288
rect 153 286 155 288
rect 149 284 155 286
rect 180 288 187 290
rect 180 286 182 288
rect 184 286 187 288
rect 133 281 138 284
rect 66 278 75 280
rect 15 267 23 273
rect 25 271 33 273
rect 25 269 28 271
rect 30 269 33 271
rect 25 267 33 269
rect 35 267 42 273
rect 55 276 62 278
rect 55 274 57 276
rect 59 274 62 276
rect 55 272 62 274
rect 57 269 62 272
rect 64 269 75 278
rect 77 269 82 280
rect 84 278 91 280
rect 84 276 87 278
rect 89 276 91 278
rect 109 279 118 281
rect 109 277 111 279
rect 113 277 118 279
rect 109 276 118 277
rect 84 274 91 276
rect 84 269 89 274
rect 97 273 102 276
rect 95 271 102 273
rect 95 269 97 271
rect 99 269 102 271
rect 95 267 102 269
rect 104 272 118 276
rect 120 276 128 281
rect 120 274 123 276
rect 125 274 128 276
rect 120 272 128 274
rect 130 278 138 281
rect 130 276 133 278
rect 135 276 138 278
rect 130 272 138 276
rect 140 272 145 284
rect 147 272 155 284
rect 180 280 187 286
rect 263 288 269 290
rect 263 286 265 288
rect 267 286 269 288
rect 263 284 269 286
rect 298 288 305 290
rect 298 286 301 288
rect 303 286 305 288
rect 247 281 252 284
rect 180 278 189 280
rect 169 276 176 278
rect 169 274 171 276
rect 173 274 176 276
rect 169 272 176 274
rect 104 267 109 272
rect 171 269 176 272
rect 178 269 189 278
rect 191 269 196 280
rect 198 278 205 280
rect 198 276 201 278
rect 203 276 205 278
rect 223 279 232 281
rect 223 277 225 279
rect 227 277 232 279
rect 223 276 232 277
rect 198 274 205 276
rect 198 269 203 274
rect 211 273 216 276
rect 209 271 216 273
rect 209 269 211 271
rect 213 269 216 271
rect 209 267 216 269
rect 218 272 232 276
rect 234 276 242 281
rect 234 274 237 276
rect 239 274 242 276
rect 234 272 242 274
rect 244 278 252 281
rect 244 276 247 278
rect 249 276 252 278
rect 244 272 252 276
rect 254 272 259 284
rect 261 272 269 284
rect 298 280 305 286
rect 280 278 287 280
rect 280 276 282 278
rect 284 276 287 278
rect 280 274 287 276
rect 218 267 223 272
rect 282 269 287 274
rect 289 269 294 280
rect 296 278 305 280
rect 333 279 339 281
rect 296 269 307 278
rect 309 276 316 278
rect 309 274 312 276
rect 314 274 316 276
rect 309 272 316 274
rect 322 277 329 279
rect 322 275 324 277
rect 326 275 329 277
rect 322 273 329 275
rect 331 277 339 279
rect 331 275 334 277
rect 336 275 339 277
rect 331 273 339 275
rect 341 273 346 281
rect 348 279 356 281
rect 348 277 351 279
rect 353 277 356 279
rect 348 273 356 277
rect 358 273 363 281
rect 365 279 373 281
rect 365 277 368 279
rect 370 277 373 279
rect 365 273 373 277
rect 309 269 314 272
rect 368 272 373 273
rect 375 278 380 281
rect 391 278 396 281
rect 375 276 382 278
rect 375 274 378 276
rect 380 274 382 276
rect 375 272 382 274
rect 389 276 396 278
rect 389 274 391 276
rect 393 274 396 276
rect 389 272 396 274
rect 398 279 406 281
rect 398 277 401 279
rect 403 277 406 279
rect 398 273 406 277
rect 408 273 413 281
rect 415 279 423 281
rect 415 277 418 279
rect 420 277 423 279
rect 415 273 423 277
rect 425 273 430 281
rect 432 279 438 281
rect 432 277 440 279
rect 432 275 435 277
rect 437 275 440 277
rect 432 273 440 275
rect 442 277 449 279
rect 458 278 463 281
rect 442 275 445 277
rect 447 275 449 277
rect 442 273 449 275
rect 456 276 463 278
rect 456 274 458 276
rect 460 274 463 276
rect 398 272 403 273
rect 456 272 463 274
rect 465 279 473 281
rect 465 277 468 279
rect 470 277 473 279
rect 465 273 473 277
rect 475 273 480 281
rect 482 279 490 281
rect 482 277 485 279
rect 487 277 490 279
rect 482 273 490 277
rect 492 273 497 281
rect 499 279 505 281
rect 564 288 570 290
rect 564 286 566 288
rect 568 286 570 288
rect 533 284 539 286
rect 533 282 535 284
rect 537 282 539 284
rect 499 277 507 279
rect 499 275 502 277
rect 504 275 507 277
rect 499 273 507 275
rect 509 277 516 279
rect 509 275 512 277
rect 514 275 516 277
rect 533 280 539 282
rect 552 284 558 286
rect 552 282 554 284
rect 556 282 558 284
rect 552 280 558 282
rect 533 276 537 280
rect 509 273 516 275
rect 524 273 529 276
rect 465 272 470 273
rect 522 271 529 273
rect 522 269 524 271
rect 526 269 529 271
rect 522 267 529 269
rect 531 273 537 276
rect 553 273 558 280
rect 531 267 539 273
rect 541 271 549 273
rect 541 269 544 271
rect 546 269 549 271
rect 541 267 549 269
rect 551 267 558 273
rect 564 284 570 286
rect 564 272 572 284
rect 574 272 579 284
rect 581 281 586 284
rect 581 278 589 281
rect 581 276 584 278
rect 586 276 589 278
rect 581 272 589 276
rect 591 276 599 281
rect 591 274 594 276
rect 596 274 599 276
rect 591 272 599 274
rect 601 279 610 281
rect 601 277 606 279
rect 608 277 610 279
rect 601 276 610 277
rect 601 272 615 276
rect 610 267 615 272
rect 617 273 622 276
rect 617 271 624 273
rect 617 269 620 271
rect 622 269 624 271
rect 617 267 624 269
rect 6 173 13 175
rect 6 171 8 173
rect 10 171 13 173
rect 6 169 13 171
rect 8 166 13 169
rect 15 169 23 175
rect 25 173 33 175
rect 25 171 28 173
rect 30 171 33 173
rect 25 169 33 171
rect 35 169 42 175
rect 95 173 102 175
rect 57 170 62 173
rect 15 166 21 169
rect 17 162 21 166
rect 37 162 42 169
rect 55 168 62 170
rect 55 166 57 168
rect 59 166 62 168
rect 55 164 62 166
rect 64 164 75 173
rect 17 160 23 162
rect 17 158 19 160
rect 21 158 23 160
rect 17 156 23 158
rect 36 160 42 162
rect 66 162 75 164
rect 77 162 82 173
rect 84 168 89 173
rect 95 171 97 173
rect 99 171 102 173
rect 95 169 102 171
rect 84 166 91 168
rect 97 166 102 169
rect 104 170 109 175
rect 209 173 216 175
rect 171 170 176 173
rect 104 166 118 170
rect 84 164 87 166
rect 89 164 91 166
rect 84 162 91 164
rect 109 165 118 166
rect 109 163 111 165
rect 113 163 118 165
rect 36 158 38 160
rect 40 158 42 160
rect 36 156 42 158
rect 66 156 73 162
rect 109 161 118 163
rect 120 168 128 170
rect 120 166 123 168
rect 125 166 128 168
rect 120 161 128 166
rect 130 166 138 170
rect 130 164 133 166
rect 135 164 138 166
rect 130 161 138 164
rect 66 154 68 156
rect 70 154 73 156
rect 66 152 73 154
rect 133 158 138 161
rect 140 158 145 170
rect 147 158 155 170
rect 169 168 176 170
rect 169 166 171 168
rect 173 166 176 168
rect 169 164 176 166
rect 178 164 189 173
rect 180 162 189 164
rect 191 162 196 173
rect 198 168 203 173
rect 209 171 211 173
rect 213 171 216 173
rect 209 169 216 171
rect 198 166 205 168
rect 211 166 216 169
rect 218 170 223 175
rect 218 166 232 170
rect 198 164 201 166
rect 203 164 205 166
rect 198 162 205 164
rect 223 165 232 166
rect 223 163 225 165
rect 227 163 232 165
rect 149 156 155 158
rect 149 154 151 156
rect 153 154 155 156
rect 149 152 155 154
rect 180 156 187 162
rect 223 161 232 163
rect 234 168 242 170
rect 234 166 237 168
rect 239 166 242 168
rect 234 161 242 166
rect 244 166 252 170
rect 244 164 247 166
rect 249 164 252 166
rect 244 161 252 164
rect 180 154 182 156
rect 184 154 187 156
rect 180 152 187 154
rect 247 158 252 161
rect 254 158 259 170
rect 261 158 269 170
rect 282 168 287 173
rect 280 166 287 168
rect 280 164 282 166
rect 284 164 287 166
rect 280 162 287 164
rect 289 162 294 173
rect 296 164 307 173
rect 309 170 314 173
rect 309 168 316 170
rect 368 169 373 170
rect 309 166 312 168
rect 314 166 316 168
rect 309 164 316 166
rect 322 167 329 169
rect 322 165 324 167
rect 326 165 329 167
rect 296 162 305 164
rect 263 156 269 158
rect 263 154 265 156
rect 267 154 269 156
rect 263 152 269 154
rect 298 156 305 162
rect 322 163 329 165
rect 331 167 339 169
rect 331 165 334 167
rect 336 165 339 167
rect 331 163 339 165
rect 298 154 301 156
rect 303 154 305 156
rect 298 152 305 154
rect 333 161 339 163
rect 341 161 346 169
rect 348 165 356 169
rect 348 163 351 165
rect 353 163 356 165
rect 348 161 356 163
rect 358 161 363 169
rect 365 165 373 169
rect 365 163 368 165
rect 370 163 373 165
rect 365 161 373 163
rect 375 168 382 170
rect 375 166 378 168
rect 380 166 382 168
rect 375 164 382 166
rect 389 168 396 170
rect 389 166 391 168
rect 393 166 396 168
rect 389 164 396 166
rect 375 161 380 164
rect 391 161 396 164
rect 398 169 403 170
rect 398 165 406 169
rect 398 163 401 165
rect 403 163 406 165
rect 398 161 406 163
rect 408 161 413 169
rect 415 165 423 169
rect 415 163 418 165
rect 420 163 423 165
rect 415 161 423 163
rect 425 161 430 169
rect 432 167 440 169
rect 432 165 435 167
rect 437 165 440 167
rect 432 163 440 165
rect 442 167 449 169
rect 442 165 445 167
rect 447 165 449 167
rect 442 163 449 165
rect 456 168 463 170
rect 456 166 458 168
rect 460 166 463 168
rect 456 164 463 166
rect 432 161 438 163
rect 458 161 463 164
rect 465 169 470 170
rect 522 173 529 175
rect 522 171 524 173
rect 526 171 529 173
rect 522 169 529 171
rect 465 165 473 169
rect 465 163 468 165
rect 470 163 473 165
rect 465 161 473 163
rect 475 161 480 169
rect 482 165 490 169
rect 482 163 485 165
rect 487 163 490 165
rect 482 161 490 163
rect 492 161 497 169
rect 499 167 507 169
rect 499 165 502 167
rect 504 165 507 167
rect 499 163 507 165
rect 509 167 516 169
rect 509 165 512 167
rect 514 165 516 167
rect 524 166 529 169
rect 531 169 539 175
rect 541 173 549 175
rect 541 171 544 173
rect 546 171 549 173
rect 541 169 549 171
rect 551 169 558 175
rect 610 170 615 175
rect 531 166 537 169
rect 509 163 516 165
rect 499 161 505 163
rect 533 162 537 166
rect 553 162 558 169
rect 533 160 539 162
rect 533 158 535 160
rect 537 158 539 160
rect 533 156 539 158
rect 552 160 558 162
rect 552 158 554 160
rect 556 158 558 160
rect 552 156 558 158
rect 564 158 572 170
rect 574 158 579 170
rect 581 166 589 170
rect 581 164 584 166
rect 586 164 589 166
rect 581 161 589 164
rect 591 168 599 170
rect 591 166 594 168
rect 596 166 599 168
rect 591 161 599 166
rect 601 166 615 170
rect 617 173 624 175
rect 617 171 620 173
rect 622 171 624 173
rect 617 169 624 171
rect 617 166 622 169
rect 601 165 610 166
rect 601 163 606 165
rect 608 163 610 165
rect 601 161 610 163
rect 581 158 586 161
rect 564 156 570 158
rect 564 154 566 156
rect 568 154 570 156
rect 564 152 570 154
rect 17 140 23 142
rect 17 138 19 140
rect 21 138 23 140
rect 17 136 23 138
rect 36 140 42 142
rect 66 144 73 146
rect 66 142 68 144
rect 70 142 73 144
rect 36 138 38 140
rect 40 138 42 140
rect 36 136 42 138
rect 17 132 21 136
rect 8 129 13 132
rect 6 127 13 129
rect 6 125 8 127
rect 10 125 13 127
rect 6 123 13 125
rect 15 129 21 132
rect 37 129 42 136
rect 66 136 73 142
rect 149 144 155 146
rect 149 142 151 144
rect 153 142 155 144
rect 149 140 155 142
rect 180 144 187 146
rect 180 142 182 144
rect 184 142 187 144
rect 133 137 138 140
rect 66 134 75 136
rect 15 123 23 129
rect 25 127 33 129
rect 25 125 28 127
rect 30 125 33 127
rect 25 123 33 125
rect 35 123 42 129
rect 55 132 62 134
rect 55 130 57 132
rect 59 130 62 132
rect 55 128 62 130
rect 57 125 62 128
rect 64 125 75 134
rect 77 125 82 136
rect 84 134 91 136
rect 84 132 87 134
rect 89 132 91 134
rect 109 135 118 137
rect 109 133 111 135
rect 113 133 118 135
rect 109 132 118 133
rect 84 130 91 132
rect 84 125 89 130
rect 97 129 102 132
rect 95 127 102 129
rect 95 125 97 127
rect 99 125 102 127
rect 95 123 102 125
rect 104 128 118 132
rect 120 132 128 137
rect 120 130 123 132
rect 125 130 128 132
rect 120 128 128 130
rect 130 134 138 137
rect 130 132 133 134
rect 135 132 138 134
rect 130 128 138 132
rect 140 128 145 140
rect 147 128 155 140
rect 180 136 187 142
rect 263 144 269 146
rect 263 142 265 144
rect 267 142 269 144
rect 263 140 269 142
rect 298 144 305 146
rect 298 142 301 144
rect 303 142 305 144
rect 247 137 252 140
rect 180 134 189 136
rect 169 132 176 134
rect 169 130 171 132
rect 173 130 176 132
rect 169 128 176 130
rect 104 123 109 128
rect 171 125 176 128
rect 178 125 189 134
rect 191 125 196 136
rect 198 134 205 136
rect 198 132 201 134
rect 203 132 205 134
rect 223 135 232 137
rect 223 133 225 135
rect 227 133 232 135
rect 223 132 232 133
rect 198 130 205 132
rect 198 125 203 130
rect 211 129 216 132
rect 209 127 216 129
rect 209 125 211 127
rect 213 125 216 127
rect 209 123 216 125
rect 218 128 232 132
rect 234 132 242 137
rect 234 130 237 132
rect 239 130 242 132
rect 234 128 242 130
rect 244 134 252 137
rect 244 132 247 134
rect 249 132 252 134
rect 244 128 252 132
rect 254 128 259 140
rect 261 128 269 140
rect 298 136 305 142
rect 280 134 287 136
rect 280 132 282 134
rect 284 132 287 134
rect 280 130 287 132
rect 218 123 223 128
rect 282 125 287 130
rect 289 125 294 136
rect 296 134 305 136
rect 333 135 339 137
rect 296 125 307 134
rect 309 132 316 134
rect 309 130 312 132
rect 314 130 316 132
rect 309 128 316 130
rect 322 133 329 135
rect 322 131 324 133
rect 326 131 329 133
rect 322 129 329 131
rect 331 133 339 135
rect 331 131 334 133
rect 336 131 339 133
rect 331 129 339 131
rect 341 129 346 137
rect 348 135 356 137
rect 348 133 351 135
rect 353 133 356 135
rect 348 129 356 133
rect 358 129 363 137
rect 365 135 373 137
rect 365 133 368 135
rect 370 133 373 135
rect 365 129 373 133
rect 309 125 314 128
rect 368 128 373 129
rect 375 134 380 137
rect 391 134 396 137
rect 375 132 382 134
rect 375 130 378 132
rect 380 130 382 132
rect 375 128 382 130
rect 389 132 396 134
rect 389 130 391 132
rect 393 130 396 132
rect 389 128 396 130
rect 398 135 406 137
rect 398 133 401 135
rect 403 133 406 135
rect 398 129 406 133
rect 408 129 413 137
rect 415 135 423 137
rect 415 133 418 135
rect 420 133 423 135
rect 415 129 423 133
rect 425 129 430 137
rect 432 135 438 137
rect 432 133 440 135
rect 432 131 435 133
rect 437 131 440 133
rect 432 129 440 131
rect 442 133 449 135
rect 458 134 463 137
rect 442 131 445 133
rect 447 131 449 133
rect 442 129 449 131
rect 456 132 463 134
rect 456 130 458 132
rect 460 130 463 132
rect 398 128 403 129
rect 456 128 463 130
rect 465 135 473 137
rect 465 133 468 135
rect 470 133 473 135
rect 465 129 473 133
rect 475 129 480 137
rect 482 135 490 137
rect 482 133 485 135
rect 487 133 490 135
rect 482 129 490 133
rect 492 129 497 137
rect 499 135 505 137
rect 564 144 570 146
rect 564 142 566 144
rect 568 142 570 144
rect 533 140 539 142
rect 533 138 535 140
rect 537 138 539 140
rect 499 133 507 135
rect 499 131 502 133
rect 504 131 507 133
rect 499 129 507 131
rect 509 133 516 135
rect 509 131 512 133
rect 514 131 516 133
rect 533 136 539 138
rect 552 140 558 142
rect 552 138 554 140
rect 556 138 558 140
rect 552 136 558 138
rect 533 132 537 136
rect 509 129 516 131
rect 524 129 529 132
rect 465 128 470 129
rect 522 127 529 129
rect 522 125 524 127
rect 526 125 529 127
rect 522 123 529 125
rect 531 129 537 132
rect 553 129 558 136
rect 531 123 539 129
rect 541 127 549 129
rect 541 125 544 127
rect 546 125 549 127
rect 541 123 549 125
rect 551 123 558 129
rect 564 140 570 142
rect 564 128 572 140
rect 574 128 579 140
rect 581 137 586 140
rect 581 134 589 137
rect 581 132 584 134
rect 586 132 589 134
rect 581 128 589 132
rect 591 132 599 137
rect 591 130 594 132
rect 596 130 599 132
rect 591 128 599 130
rect 601 135 610 137
rect 601 133 606 135
rect 608 133 610 135
rect 601 132 610 133
rect 601 128 615 132
rect 610 123 615 128
rect 617 129 622 132
rect 617 127 624 129
rect 617 125 620 127
rect 622 125 624 127
rect 617 123 624 125
rect 6 29 13 31
rect 6 27 8 29
rect 10 27 13 29
rect 6 25 13 27
rect 8 22 13 25
rect 15 25 23 31
rect 25 29 33 31
rect 25 27 28 29
rect 30 27 33 29
rect 25 25 33 27
rect 35 25 42 31
rect 95 29 102 31
rect 57 26 62 29
rect 15 22 21 25
rect 17 18 21 22
rect 37 18 42 25
rect 55 24 62 26
rect 55 22 57 24
rect 59 22 62 24
rect 55 20 62 22
rect 64 20 75 29
rect 17 16 23 18
rect 17 14 19 16
rect 21 14 23 16
rect 17 12 23 14
rect 36 16 42 18
rect 66 18 75 20
rect 77 18 82 29
rect 84 24 89 29
rect 95 27 97 29
rect 99 27 102 29
rect 95 25 102 27
rect 84 22 91 24
rect 97 22 102 25
rect 104 26 109 31
rect 209 29 216 31
rect 171 26 176 29
rect 104 22 118 26
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 109 21 118 22
rect 109 19 111 21
rect 113 19 118 21
rect 36 14 38 16
rect 40 14 42 16
rect 36 12 42 14
rect 66 12 73 18
rect 109 17 118 19
rect 120 24 128 26
rect 120 22 123 24
rect 125 22 128 24
rect 120 17 128 22
rect 130 22 138 26
rect 130 20 133 22
rect 135 20 138 22
rect 130 17 138 20
rect 66 10 68 12
rect 70 10 73 12
rect 66 8 73 10
rect 133 14 138 17
rect 140 14 145 26
rect 147 14 155 26
rect 169 24 176 26
rect 169 22 171 24
rect 173 22 176 24
rect 169 20 176 22
rect 178 20 189 29
rect 180 18 189 20
rect 191 18 196 29
rect 198 24 203 29
rect 209 27 211 29
rect 213 27 216 29
rect 209 25 216 27
rect 198 22 205 24
rect 211 22 216 25
rect 218 26 223 31
rect 218 22 232 26
rect 198 20 201 22
rect 203 20 205 22
rect 198 18 205 20
rect 223 21 232 22
rect 223 19 225 21
rect 227 19 232 21
rect 149 12 155 14
rect 149 10 151 12
rect 153 10 155 12
rect 149 8 155 10
rect 180 12 187 18
rect 223 17 232 19
rect 234 24 242 26
rect 234 22 237 24
rect 239 22 242 24
rect 234 17 242 22
rect 244 22 252 26
rect 244 20 247 22
rect 249 20 252 22
rect 244 17 252 20
rect 180 10 182 12
rect 184 10 187 12
rect 180 8 187 10
rect 247 14 252 17
rect 254 14 259 26
rect 261 14 269 26
rect 282 24 287 29
rect 280 22 287 24
rect 280 20 282 22
rect 284 20 287 22
rect 280 18 287 20
rect 289 18 294 29
rect 296 20 307 29
rect 309 26 314 29
rect 309 24 316 26
rect 368 25 373 26
rect 309 22 312 24
rect 314 22 316 24
rect 309 20 316 22
rect 322 23 329 25
rect 322 21 324 23
rect 326 21 329 23
rect 296 18 305 20
rect 263 12 269 14
rect 263 10 265 12
rect 267 10 269 12
rect 263 8 269 10
rect 298 12 305 18
rect 322 19 329 21
rect 331 23 339 25
rect 331 21 334 23
rect 336 21 339 23
rect 331 19 339 21
rect 298 10 301 12
rect 303 10 305 12
rect 298 8 305 10
rect 333 17 339 19
rect 341 17 346 25
rect 348 21 356 25
rect 348 19 351 21
rect 353 19 356 21
rect 348 17 356 19
rect 358 17 363 25
rect 365 21 373 25
rect 365 19 368 21
rect 370 19 373 21
rect 365 17 373 19
rect 375 24 382 26
rect 375 22 378 24
rect 380 22 382 24
rect 375 20 382 22
rect 389 24 396 26
rect 389 22 391 24
rect 393 22 396 24
rect 389 20 396 22
rect 375 17 380 20
rect 391 17 396 20
rect 398 25 403 26
rect 398 21 406 25
rect 398 19 401 21
rect 403 19 406 21
rect 398 17 406 19
rect 408 17 413 25
rect 415 21 423 25
rect 415 19 418 21
rect 420 19 423 21
rect 415 17 423 19
rect 425 17 430 25
rect 432 23 440 25
rect 432 21 435 23
rect 437 21 440 23
rect 432 19 440 21
rect 442 23 449 25
rect 442 21 445 23
rect 447 21 449 23
rect 442 19 449 21
rect 456 24 463 26
rect 456 22 458 24
rect 460 22 463 24
rect 456 20 463 22
rect 432 17 438 19
rect 458 17 463 20
rect 465 25 470 26
rect 522 29 529 31
rect 522 27 524 29
rect 526 27 529 29
rect 522 25 529 27
rect 465 21 473 25
rect 465 19 468 21
rect 470 19 473 21
rect 465 17 473 19
rect 475 17 480 25
rect 482 21 490 25
rect 482 19 485 21
rect 487 19 490 21
rect 482 17 490 19
rect 492 17 497 25
rect 499 23 507 25
rect 499 21 502 23
rect 504 21 507 23
rect 499 19 507 21
rect 509 23 516 25
rect 509 21 512 23
rect 514 21 516 23
rect 524 22 529 25
rect 531 25 539 31
rect 541 29 549 31
rect 541 27 544 29
rect 546 27 549 29
rect 541 25 549 27
rect 551 25 558 31
rect 610 26 615 31
rect 531 22 537 25
rect 509 19 516 21
rect 499 17 505 19
rect 533 18 537 22
rect 553 18 558 25
rect 533 16 539 18
rect 533 14 535 16
rect 537 14 539 16
rect 533 12 539 14
rect 552 16 558 18
rect 552 14 554 16
rect 556 14 558 16
rect 552 12 558 14
rect 564 14 572 26
rect 574 14 579 26
rect 581 22 589 26
rect 581 20 584 22
rect 586 20 589 22
rect 581 17 589 20
rect 591 24 599 26
rect 591 22 594 24
rect 596 22 599 24
rect 591 17 599 22
rect 601 22 615 26
rect 617 29 624 31
rect 617 27 620 29
rect 622 27 624 29
rect 617 25 624 27
rect 617 22 622 25
rect 601 21 610 22
rect 601 19 606 21
rect 608 19 610 21
rect 601 17 610 19
rect 581 14 586 17
rect 564 12 570 14
rect 564 10 566 12
rect 568 10 570 12
rect 564 8 570 10
<< pdif >>
rect 8 250 13 255
rect 6 248 13 250
rect 6 246 8 248
rect 10 246 13 248
rect 6 241 13 246
rect 6 239 8 241
rect 10 239 13 241
rect 6 237 13 239
rect 15 248 23 255
rect 55 252 62 254
rect 55 250 57 252
rect 59 250 62 252
rect 15 237 26 248
rect 17 231 26 237
rect 17 229 19 231
rect 21 229 26 231
rect 17 227 26 229
rect 28 227 33 248
rect 35 240 40 248
rect 55 245 62 250
rect 55 243 57 245
rect 59 243 62 245
rect 55 241 62 243
rect 35 238 42 240
rect 35 236 38 238
rect 40 236 42 238
rect 57 236 62 241
rect 64 247 70 254
rect 103 252 110 254
rect 103 250 105 252
rect 107 250 110 252
rect 103 248 110 250
rect 64 240 72 247
rect 64 238 67 240
rect 69 238 72 240
rect 64 236 72 238
rect 35 234 42 236
rect 35 227 40 234
rect 66 234 72 236
rect 74 245 82 247
rect 74 243 77 245
rect 79 243 82 245
rect 74 238 82 243
rect 74 236 77 238
rect 79 236 82 238
rect 74 234 82 236
rect 84 238 91 247
rect 84 236 87 238
rect 89 236 91 238
rect 84 234 91 236
rect 105 227 110 248
rect 112 238 126 254
rect 112 236 115 238
rect 117 236 126 238
rect 128 252 136 254
rect 128 250 131 252
rect 133 250 136 252
rect 128 245 136 250
rect 128 243 131 245
rect 133 243 136 245
rect 128 236 136 243
rect 138 245 146 254
rect 138 243 141 245
rect 143 243 146 245
rect 138 236 146 243
rect 112 231 124 236
rect 112 229 115 231
rect 117 229 124 231
rect 112 227 124 229
rect 141 227 146 236
rect 148 239 153 254
rect 169 252 176 254
rect 169 250 171 252
rect 173 250 176 252
rect 169 245 176 250
rect 169 243 171 245
rect 173 243 176 245
rect 169 241 176 243
rect 148 237 155 239
rect 148 235 151 237
rect 153 235 155 237
rect 171 236 176 241
rect 178 247 184 254
rect 217 252 224 254
rect 217 250 219 252
rect 221 250 224 252
rect 217 248 224 250
rect 178 240 186 247
rect 178 238 181 240
rect 183 238 186 240
rect 178 236 186 238
rect 148 233 155 235
rect 148 227 153 233
rect 180 234 186 236
rect 188 245 196 247
rect 188 243 191 245
rect 193 243 196 245
rect 188 238 196 243
rect 188 236 191 238
rect 193 236 196 238
rect 188 234 196 236
rect 198 238 205 247
rect 198 236 201 238
rect 203 236 205 238
rect 198 234 205 236
rect 219 227 224 248
rect 226 238 240 254
rect 226 236 229 238
rect 231 236 240 238
rect 242 252 250 254
rect 242 250 245 252
rect 247 250 250 252
rect 242 245 250 250
rect 242 243 245 245
rect 247 243 250 245
rect 242 236 250 243
rect 252 245 260 254
rect 252 243 255 245
rect 257 243 260 245
rect 252 236 260 243
rect 226 231 238 236
rect 226 229 229 231
rect 231 229 238 231
rect 226 227 238 229
rect 255 227 260 236
rect 262 239 267 254
rect 301 247 307 254
rect 262 237 269 239
rect 262 235 265 237
rect 267 235 269 237
rect 262 233 269 235
rect 280 238 287 247
rect 280 236 282 238
rect 284 236 287 238
rect 280 234 287 236
rect 289 245 297 247
rect 289 243 292 245
rect 294 243 297 245
rect 289 238 297 243
rect 289 236 292 238
rect 294 236 297 238
rect 289 234 297 236
rect 299 240 307 247
rect 299 238 302 240
rect 304 238 307 240
rect 299 236 307 238
rect 309 252 316 254
rect 309 250 312 252
rect 314 250 316 252
rect 309 245 316 250
rect 322 253 329 255
rect 322 251 324 253
rect 326 251 329 253
rect 322 249 329 251
rect 324 247 329 249
rect 331 247 337 255
rect 309 243 312 245
rect 314 243 316 245
rect 309 241 316 243
rect 333 243 337 247
rect 368 243 373 245
rect 309 236 314 241
rect 333 239 339 243
rect 299 234 305 236
rect 262 227 267 233
rect 332 231 339 239
rect 332 229 334 231
rect 336 229 339 231
rect 332 227 339 229
rect 341 227 346 243
rect 348 241 356 243
rect 348 239 351 241
rect 353 239 356 241
rect 348 227 356 239
rect 358 227 363 243
rect 365 231 373 243
rect 365 229 368 231
rect 370 229 373 231
rect 365 227 373 229
rect 375 240 380 245
rect 391 240 396 245
rect 375 238 382 240
rect 375 236 378 238
rect 380 236 382 238
rect 375 234 382 236
rect 389 238 396 240
rect 389 236 391 238
rect 393 236 396 238
rect 389 234 396 236
rect 375 227 380 234
rect 391 227 396 234
rect 398 243 403 245
rect 434 247 440 255
rect 442 253 449 255
rect 442 251 445 253
rect 447 251 449 253
rect 442 249 449 251
rect 442 247 447 249
rect 434 243 438 247
rect 398 231 406 243
rect 398 229 401 231
rect 403 229 406 231
rect 398 227 406 229
rect 408 227 413 243
rect 415 241 423 243
rect 415 239 418 241
rect 420 239 423 241
rect 415 227 423 239
rect 425 227 430 243
rect 432 239 438 243
rect 458 240 463 245
rect 432 231 439 239
rect 456 238 463 240
rect 456 236 458 238
rect 460 236 463 238
rect 456 234 463 236
rect 432 229 435 231
rect 437 229 439 231
rect 432 227 439 229
rect 458 227 463 234
rect 465 243 470 245
rect 501 247 507 255
rect 509 253 516 255
rect 509 251 512 253
rect 514 251 516 253
rect 509 249 516 251
rect 524 250 529 255
rect 509 247 514 249
rect 522 248 529 250
rect 501 243 505 247
rect 465 231 473 243
rect 465 229 468 231
rect 470 229 473 231
rect 465 227 473 229
rect 475 227 480 243
rect 482 241 490 243
rect 482 239 485 241
rect 487 239 490 241
rect 482 227 490 239
rect 492 227 497 243
rect 499 239 505 243
rect 522 246 524 248
rect 526 246 529 248
rect 499 231 506 239
rect 522 241 529 246
rect 522 239 524 241
rect 526 239 529 241
rect 522 237 529 239
rect 531 248 539 255
rect 531 237 542 248
rect 499 229 502 231
rect 504 229 506 231
rect 533 231 542 237
rect 499 227 506 229
rect 533 229 535 231
rect 537 229 542 231
rect 533 227 542 229
rect 544 227 549 248
rect 551 240 556 248
rect 551 238 558 240
rect 566 239 571 254
rect 551 236 554 238
rect 556 236 558 238
rect 551 234 558 236
rect 564 237 571 239
rect 564 235 566 237
rect 568 235 571 237
rect 551 227 556 234
rect 564 233 571 235
rect 566 227 571 233
rect 573 245 581 254
rect 573 243 576 245
rect 578 243 581 245
rect 573 236 581 243
rect 583 252 591 254
rect 583 250 586 252
rect 588 250 591 252
rect 583 245 591 250
rect 583 243 586 245
rect 588 243 591 245
rect 583 236 591 243
rect 593 238 607 254
rect 593 236 602 238
rect 604 236 607 238
rect 573 227 578 236
rect 595 231 607 236
rect 595 229 602 231
rect 604 229 607 231
rect 595 227 607 229
rect 609 252 616 254
rect 609 250 612 252
rect 614 250 616 252
rect 609 248 616 250
rect 609 227 614 248
rect 17 213 26 215
rect 17 211 19 213
rect 21 211 26 213
rect 17 205 26 211
rect 6 203 13 205
rect 6 201 8 203
rect 10 201 13 203
rect 6 196 13 201
rect 6 194 8 196
rect 10 194 13 196
rect 6 192 13 194
rect 8 187 13 192
rect 15 194 26 205
rect 28 194 33 215
rect 35 208 40 215
rect 35 206 42 208
rect 66 206 72 208
rect 35 204 38 206
rect 40 204 42 206
rect 35 202 42 204
rect 35 194 40 202
rect 57 201 62 206
rect 55 199 62 201
rect 55 197 57 199
rect 59 197 62 199
rect 15 187 23 194
rect 55 192 62 197
rect 55 190 57 192
rect 59 190 62 192
rect 55 188 62 190
rect 64 204 72 206
rect 64 202 67 204
rect 69 202 72 204
rect 64 195 72 202
rect 74 206 82 208
rect 74 204 77 206
rect 79 204 82 206
rect 74 199 82 204
rect 74 197 77 199
rect 79 197 82 199
rect 74 195 82 197
rect 84 206 91 208
rect 84 204 87 206
rect 89 204 91 206
rect 84 195 91 204
rect 64 188 70 195
rect 105 194 110 215
rect 103 192 110 194
rect 103 190 105 192
rect 107 190 110 192
rect 103 188 110 190
rect 112 213 124 215
rect 112 211 115 213
rect 117 211 124 213
rect 112 206 124 211
rect 141 206 146 215
rect 112 204 115 206
rect 117 204 126 206
rect 112 188 126 204
rect 128 199 136 206
rect 128 197 131 199
rect 133 197 136 199
rect 128 192 136 197
rect 128 190 131 192
rect 133 190 136 192
rect 128 188 136 190
rect 138 199 146 206
rect 138 197 141 199
rect 143 197 146 199
rect 138 188 146 197
rect 148 209 153 215
rect 148 207 155 209
rect 148 205 151 207
rect 153 205 155 207
rect 180 206 186 208
rect 148 203 155 205
rect 148 188 153 203
rect 171 201 176 206
rect 169 199 176 201
rect 169 197 171 199
rect 173 197 176 199
rect 169 192 176 197
rect 169 190 171 192
rect 173 190 176 192
rect 169 188 176 190
rect 178 204 186 206
rect 178 202 181 204
rect 183 202 186 204
rect 178 195 186 202
rect 188 206 196 208
rect 188 204 191 206
rect 193 204 196 206
rect 188 199 196 204
rect 188 197 191 199
rect 193 197 196 199
rect 188 195 196 197
rect 198 206 205 208
rect 198 204 201 206
rect 203 204 205 206
rect 198 195 205 204
rect 178 188 184 195
rect 219 194 224 215
rect 217 192 224 194
rect 217 190 219 192
rect 221 190 224 192
rect 217 188 224 190
rect 226 213 238 215
rect 226 211 229 213
rect 231 211 238 213
rect 226 206 238 211
rect 255 206 260 215
rect 226 204 229 206
rect 231 204 240 206
rect 226 188 240 204
rect 242 199 250 206
rect 242 197 245 199
rect 247 197 250 199
rect 242 192 250 197
rect 242 190 245 192
rect 247 190 250 192
rect 242 188 250 190
rect 252 199 260 206
rect 252 197 255 199
rect 257 197 260 199
rect 252 188 260 197
rect 262 209 267 215
rect 262 207 269 209
rect 332 213 339 215
rect 332 211 334 213
rect 336 211 339 213
rect 262 205 265 207
rect 267 205 269 207
rect 262 203 269 205
rect 280 206 287 208
rect 280 204 282 206
rect 284 204 287 206
rect 262 188 267 203
rect 280 195 287 204
rect 289 206 297 208
rect 289 204 292 206
rect 294 204 297 206
rect 289 199 297 204
rect 289 197 292 199
rect 294 197 297 199
rect 289 195 297 197
rect 299 206 305 208
rect 299 204 307 206
rect 299 202 302 204
rect 304 202 307 204
rect 299 195 307 202
rect 301 188 307 195
rect 309 201 314 206
rect 332 203 339 211
rect 309 199 316 201
rect 309 197 312 199
rect 314 197 316 199
rect 309 192 316 197
rect 333 199 339 203
rect 341 199 346 215
rect 348 203 356 215
rect 348 201 351 203
rect 353 201 356 203
rect 348 199 356 201
rect 358 199 363 215
rect 365 213 373 215
rect 365 211 368 213
rect 370 211 373 213
rect 365 199 373 211
rect 333 195 337 199
rect 324 193 329 195
rect 309 190 312 192
rect 314 190 316 192
rect 309 188 316 190
rect 322 191 329 193
rect 322 189 324 191
rect 326 189 329 191
rect 322 187 329 189
rect 331 187 337 195
rect 368 197 373 199
rect 375 208 380 215
rect 391 208 396 215
rect 375 206 382 208
rect 375 204 378 206
rect 380 204 382 206
rect 375 202 382 204
rect 389 206 396 208
rect 389 204 391 206
rect 393 204 396 206
rect 389 202 396 204
rect 375 197 380 202
rect 391 197 396 202
rect 398 213 406 215
rect 398 211 401 213
rect 403 211 406 213
rect 398 199 406 211
rect 408 199 413 215
rect 415 203 423 215
rect 415 201 418 203
rect 420 201 423 203
rect 415 199 423 201
rect 425 199 430 215
rect 432 213 439 215
rect 432 211 435 213
rect 437 211 439 213
rect 432 203 439 211
rect 458 208 463 215
rect 456 206 463 208
rect 456 204 458 206
rect 460 204 463 206
rect 432 199 438 203
rect 456 202 463 204
rect 398 197 403 199
rect 434 195 438 199
rect 458 197 463 202
rect 465 213 473 215
rect 465 211 468 213
rect 470 211 473 213
rect 465 199 473 211
rect 475 199 480 215
rect 482 203 490 215
rect 482 201 485 203
rect 487 201 490 203
rect 482 199 490 201
rect 492 199 497 215
rect 499 213 506 215
rect 499 211 502 213
rect 504 211 506 213
rect 533 213 542 215
rect 499 203 506 211
rect 533 211 535 213
rect 537 211 542 213
rect 533 205 542 211
rect 499 199 505 203
rect 465 197 470 199
rect 434 187 440 195
rect 442 193 447 195
rect 442 191 449 193
rect 442 189 445 191
rect 447 189 449 191
rect 442 187 449 189
rect 501 195 505 199
rect 522 203 529 205
rect 522 201 524 203
rect 526 201 529 203
rect 522 196 529 201
rect 501 187 507 195
rect 509 193 514 195
rect 522 194 524 196
rect 526 194 529 196
rect 509 191 516 193
rect 522 192 529 194
rect 509 189 512 191
rect 514 189 516 191
rect 509 187 516 189
rect 524 187 529 192
rect 531 194 542 205
rect 544 194 549 215
rect 551 208 556 215
rect 566 209 571 215
rect 551 206 558 208
rect 551 204 554 206
rect 556 204 558 206
rect 551 202 558 204
rect 564 207 571 209
rect 564 205 566 207
rect 568 205 571 207
rect 564 203 571 205
rect 551 194 556 202
rect 531 187 539 194
rect 566 188 571 203
rect 573 206 578 215
rect 595 213 607 215
rect 595 211 602 213
rect 604 211 607 213
rect 595 206 607 211
rect 573 199 581 206
rect 573 197 576 199
rect 578 197 581 199
rect 573 188 581 197
rect 583 199 591 206
rect 583 197 586 199
rect 588 197 591 199
rect 583 192 591 197
rect 583 190 586 192
rect 588 190 591 192
rect 583 188 591 190
rect 593 204 602 206
rect 604 204 607 206
rect 593 188 607 204
rect 609 194 614 215
rect 609 192 616 194
rect 609 190 612 192
rect 614 190 616 192
rect 609 188 616 190
rect 8 106 13 111
rect 6 104 13 106
rect 6 102 8 104
rect 10 102 13 104
rect 6 97 13 102
rect 6 95 8 97
rect 10 95 13 97
rect 6 93 13 95
rect 15 104 23 111
rect 55 108 62 110
rect 55 106 57 108
rect 59 106 62 108
rect 15 93 26 104
rect 17 87 26 93
rect 17 85 19 87
rect 21 85 26 87
rect 17 83 26 85
rect 28 83 33 104
rect 35 96 40 104
rect 55 101 62 106
rect 55 99 57 101
rect 59 99 62 101
rect 55 97 62 99
rect 35 94 42 96
rect 35 92 38 94
rect 40 92 42 94
rect 57 92 62 97
rect 64 103 70 110
rect 103 108 110 110
rect 103 106 105 108
rect 107 106 110 108
rect 103 104 110 106
rect 64 96 72 103
rect 64 94 67 96
rect 69 94 72 96
rect 64 92 72 94
rect 35 90 42 92
rect 35 83 40 90
rect 66 90 72 92
rect 74 101 82 103
rect 74 99 77 101
rect 79 99 82 101
rect 74 94 82 99
rect 74 92 77 94
rect 79 92 82 94
rect 74 90 82 92
rect 84 94 91 103
rect 84 92 87 94
rect 89 92 91 94
rect 84 90 91 92
rect 105 83 110 104
rect 112 94 126 110
rect 112 92 115 94
rect 117 92 126 94
rect 128 108 136 110
rect 128 106 131 108
rect 133 106 136 108
rect 128 101 136 106
rect 128 99 131 101
rect 133 99 136 101
rect 128 92 136 99
rect 138 101 146 110
rect 138 99 141 101
rect 143 99 146 101
rect 138 92 146 99
rect 112 87 124 92
rect 112 85 115 87
rect 117 85 124 87
rect 112 83 124 85
rect 141 83 146 92
rect 148 95 153 110
rect 169 108 176 110
rect 169 106 171 108
rect 173 106 176 108
rect 169 101 176 106
rect 169 99 171 101
rect 173 99 176 101
rect 169 97 176 99
rect 148 93 155 95
rect 148 91 151 93
rect 153 91 155 93
rect 171 92 176 97
rect 178 103 184 110
rect 217 108 224 110
rect 217 106 219 108
rect 221 106 224 108
rect 217 104 224 106
rect 178 96 186 103
rect 178 94 181 96
rect 183 94 186 96
rect 178 92 186 94
rect 148 89 155 91
rect 148 83 153 89
rect 180 90 186 92
rect 188 101 196 103
rect 188 99 191 101
rect 193 99 196 101
rect 188 94 196 99
rect 188 92 191 94
rect 193 92 196 94
rect 188 90 196 92
rect 198 94 205 103
rect 198 92 201 94
rect 203 92 205 94
rect 198 90 205 92
rect 219 83 224 104
rect 226 94 240 110
rect 226 92 229 94
rect 231 92 240 94
rect 242 108 250 110
rect 242 106 245 108
rect 247 106 250 108
rect 242 101 250 106
rect 242 99 245 101
rect 247 99 250 101
rect 242 92 250 99
rect 252 101 260 110
rect 252 99 255 101
rect 257 99 260 101
rect 252 92 260 99
rect 226 87 238 92
rect 226 85 229 87
rect 231 85 238 87
rect 226 83 238 85
rect 255 83 260 92
rect 262 95 267 110
rect 301 103 307 110
rect 262 93 269 95
rect 262 91 265 93
rect 267 91 269 93
rect 262 89 269 91
rect 280 94 287 103
rect 280 92 282 94
rect 284 92 287 94
rect 280 90 287 92
rect 289 101 297 103
rect 289 99 292 101
rect 294 99 297 101
rect 289 94 297 99
rect 289 92 292 94
rect 294 92 297 94
rect 289 90 297 92
rect 299 96 307 103
rect 299 94 302 96
rect 304 94 307 96
rect 299 92 307 94
rect 309 108 316 110
rect 309 106 312 108
rect 314 106 316 108
rect 309 101 316 106
rect 322 109 329 111
rect 322 107 324 109
rect 326 107 329 109
rect 322 105 329 107
rect 324 103 329 105
rect 331 103 337 111
rect 309 99 312 101
rect 314 99 316 101
rect 309 97 316 99
rect 333 99 337 103
rect 368 99 373 101
rect 309 92 314 97
rect 333 95 339 99
rect 299 90 305 92
rect 262 83 267 89
rect 332 87 339 95
rect 332 85 334 87
rect 336 85 339 87
rect 332 83 339 85
rect 341 83 346 99
rect 348 97 356 99
rect 348 95 351 97
rect 353 95 356 97
rect 348 83 356 95
rect 358 83 363 99
rect 365 87 373 99
rect 365 85 368 87
rect 370 85 373 87
rect 365 83 373 85
rect 375 96 380 101
rect 391 96 396 101
rect 375 94 382 96
rect 375 92 378 94
rect 380 92 382 94
rect 375 90 382 92
rect 389 94 396 96
rect 389 92 391 94
rect 393 92 396 94
rect 389 90 396 92
rect 375 83 380 90
rect 391 83 396 90
rect 398 99 403 101
rect 434 103 440 111
rect 442 109 449 111
rect 442 107 445 109
rect 447 107 449 109
rect 442 105 449 107
rect 442 103 447 105
rect 434 99 438 103
rect 398 87 406 99
rect 398 85 401 87
rect 403 85 406 87
rect 398 83 406 85
rect 408 83 413 99
rect 415 97 423 99
rect 415 95 418 97
rect 420 95 423 97
rect 415 83 423 95
rect 425 83 430 99
rect 432 95 438 99
rect 458 96 463 101
rect 432 87 439 95
rect 456 94 463 96
rect 456 92 458 94
rect 460 92 463 94
rect 456 90 463 92
rect 432 85 435 87
rect 437 85 439 87
rect 432 83 439 85
rect 458 83 463 90
rect 465 99 470 101
rect 501 103 507 111
rect 509 109 516 111
rect 509 107 512 109
rect 514 107 516 109
rect 509 105 516 107
rect 524 106 529 111
rect 509 103 514 105
rect 522 104 529 106
rect 501 99 505 103
rect 465 87 473 99
rect 465 85 468 87
rect 470 85 473 87
rect 465 83 473 85
rect 475 83 480 99
rect 482 97 490 99
rect 482 95 485 97
rect 487 95 490 97
rect 482 83 490 95
rect 492 83 497 99
rect 499 95 505 99
rect 522 102 524 104
rect 526 102 529 104
rect 499 87 506 95
rect 522 97 529 102
rect 522 95 524 97
rect 526 95 529 97
rect 522 93 529 95
rect 531 104 539 111
rect 531 93 542 104
rect 499 85 502 87
rect 504 85 506 87
rect 533 87 542 93
rect 499 83 506 85
rect 533 85 535 87
rect 537 85 542 87
rect 533 83 542 85
rect 544 83 549 104
rect 551 96 556 104
rect 551 94 558 96
rect 566 95 571 110
rect 551 92 554 94
rect 556 92 558 94
rect 551 90 558 92
rect 564 93 571 95
rect 564 91 566 93
rect 568 91 571 93
rect 551 83 556 90
rect 564 89 571 91
rect 566 83 571 89
rect 573 101 581 110
rect 573 99 576 101
rect 578 99 581 101
rect 573 92 581 99
rect 583 108 591 110
rect 583 106 586 108
rect 588 106 591 108
rect 583 101 591 106
rect 583 99 586 101
rect 588 99 591 101
rect 583 92 591 99
rect 593 94 607 110
rect 593 92 602 94
rect 604 92 607 94
rect 573 83 578 92
rect 595 87 607 92
rect 595 85 602 87
rect 604 85 607 87
rect 595 83 607 85
rect 609 108 616 110
rect 609 106 612 108
rect 614 106 616 108
rect 609 104 616 106
rect 609 83 614 104
rect 17 69 26 71
rect 17 67 19 69
rect 21 67 26 69
rect 17 61 26 67
rect 6 59 13 61
rect 6 57 8 59
rect 10 57 13 59
rect 6 52 13 57
rect 6 50 8 52
rect 10 50 13 52
rect 6 48 13 50
rect 8 43 13 48
rect 15 50 26 61
rect 28 50 33 71
rect 35 64 40 71
rect 35 62 42 64
rect 66 62 72 64
rect 35 60 38 62
rect 40 60 42 62
rect 35 58 42 60
rect 35 50 40 58
rect 57 57 62 62
rect 55 55 62 57
rect 55 53 57 55
rect 59 53 62 55
rect 15 43 23 50
rect 55 48 62 53
rect 55 46 57 48
rect 59 46 62 48
rect 55 44 62 46
rect 64 60 72 62
rect 64 58 67 60
rect 69 58 72 60
rect 64 51 72 58
rect 74 62 82 64
rect 74 60 77 62
rect 79 60 82 62
rect 74 55 82 60
rect 74 53 77 55
rect 79 53 82 55
rect 74 51 82 53
rect 84 62 91 64
rect 84 60 87 62
rect 89 60 91 62
rect 84 51 91 60
rect 64 44 70 51
rect 105 50 110 71
rect 103 48 110 50
rect 103 46 105 48
rect 107 46 110 48
rect 103 44 110 46
rect 112 69 124 71
rect 112 67 115 69
rect 117 67 124 69
rect 112 62 124 67
rect 141 62 146 71
rect 112 60 115 62
rect 117 60 126 62
rect 112 44 126 60
rect 128 55 136 62
rect 128 53 131 55
rect 133 53 136 55
rect 128 48 136 53
rect 128 46 131 48
rect 133 46 136 48
rect 128 44 136 46
rect 138 55 146 62
rect 138 53 141 55
rect 143 53 146 55
rect 138 44 146 53
rect 148 65 153 71
rect 148 63 155 65
rect 148 61 151 63
rect 153 61 155 63
rect 180 62 186 64
rect 148 59 155 61
rect 148 44 153 59
rect 171 57 176 62
rect 169 55 176 57
rect 169 53 171 55
rect 173 53 176 55
rect 169 48 176 53
rect 169 46 171 48
rect 173 46 176 48
rect 169 44 176 46
rect 178 60 186 62
rect 178 58 181 60
rect 183 58 186 60
rect 178 51 186 58
rect 188 62 196 64
rect 188 60 191 62
rect 193 60 196 62
rect 188 55 196 60
rect 188 53 191 55
rect 193 53 196 55
rect 188 51 196 53
rect 198 62 205 64
rect 198 60 201 62
rect 203 60 205 62
rect 198 51 205 60
rect 178 44 184 51
rect 219 50 224 71
rect 217 48 224 50
rect 217 46 219 48
rect 221 46 224 48
rect 217 44 224 46
rect 226 69 238 71
rect 226 67 229 69
rect 231 67 238 69
rect 226 62 238 67
rect 255 62 260 71
rect 226 60 229 62
rect 231 60 240 62
rect 226 44 240 60
rect 242 55 250 62
rect 242 53 245 55
rect 247 53 250 55
rect 242 48 250 53
rect 242 46 245 48
rect 247 46 250 48
rect 242 44 250 46
rect 252 55 260 62
rect 252 53 255 55
rect 257 53 260 55
rect 252 44 260 53
rect 262 65 267 71
rect 262 63 269 65
rect 332 69 339 71
rect 332 67 334 69
rect 336 67 339 69
rect 262 61 265 63
rect 267 61 269 63
rect 262 59 269 61
rect 280 62 287 64
rect 280 60 282 62
rect 284 60 287 62
rect 262 44 267 59
rect 280 51 287 60
rect 289 62 297 64
rect 289 60 292 62
rect 294 60 297 62
rect 289 55 297 60
rect 289 53 292 55
rect 294 53 297 55
rect 289 51 297 53
rect 299 62 305 64
rect 299 60 307 62
rect 299 58 302 60
rect 304 58 307 60
rect 299 51 307 58
rect 301 44 307 51
rect 309 57 314 62
rect 332 59 339 67
rect 309 55 316 57
rect 309 53 312 55
rect 314 53 316 55
rect 309 48 316 53
rect 333 55 339 59
rect 341 55 346 71
rect 348 59 356 71
rect 348 57 351 59
rect 353 57 356 59
rect 348 55 356 57
rect 358 55 363 71
rect 365 69 373 71
rect 365 67 368 69
rect 370 67 373 69
rect 365 55 373 67
rect 333 51 337 55
rect 324 49 329 51
rect 309 46 312 48
rect 314 46 316 48
rect 309 44 316 46
rect 322 47 329 49
rect 322 45 324 47
rect 326 45 329 47
rect 322 43 329 45
rect 331 43 337 51
rect 368 53 373 55
rect 375 64 380 71
rect 391 64 396 71
rect 375 62 382 64
rect 375 60 378 62
rect 380 60 382 62
rect 375 58 382 60
rect 389 62 396 64
rect 389 60 391 62
rect 393 60 396 62
rect 389 58 396 60
rect 375 53 380 58
rect 391 53 396 58
rect 398 69 406 71
rect 398 67 401 69
rect 403 67 406 69
rect 398 55 406 67
rect 408 55 413 71
rect 415 59 423 71
rect 415 57 418 59
rect 420 57 423 59
rect 415 55 423 57
rect 425 55 430 71
rect 432 69 439 71
rect 432 67 435 69
rect 437 67 439 69
rect 432 59 439 67
rect 458 64 463 71
rect 456 62 463 64
rect 456 60 458 62
rect 460 60 463 62
rect 432 55 438 59
rect 456 58 463 60
rect 398 53 403 55
rect 434 51 438 55
rect 458 53 463 58
rect 465 69 473 71
rect 465 67 468 69
rect 470 67 473 69
rect 465 55 473 67
rect 475 55 480 71
rect 482 59 490 71
rect 482 57 485 59
rect 487 57 490 59
rect 482 55 490 57
rect 492 55 497 71
rect 499 69 506 71
rect 499 67 502 69
rect 504 67 506 69
rect 533 69 542 71
rect 499 59 506 67
rect 533 67 535 69
rect 537 67 542 69
rect 533 61 542 67
rect 499 55 505 59
rect 465 53 470 55
rect 434 43 440 51
rect 442 49 447 51
rect 442 47 449 49
rect 442 45 445 47
rect 447 45 449 47
rect 442 43 449 45
rect 501 51 505 55
rect 522 59 529 61
rect 522 57 524 59
rect 526 57 529 59
rect 522 52 529 57
rect 501 43 507 51
rect 509 49 514 51
rect 522 50 524 52
rect 526 50 529 52
rect 509 47 516 49
rect 522 48 529 50
rect 509 45 512 47
rect 514 45 516 47
rect 509 43 516 45
rect 524 43 529 48
rect 531 50 542 61
rect 544 50 549 71
rect 551 64 556 71
rect 566 65 571 71
rect 551 62 558 64
rect 551 60 554 62
rect 556 60 558 62
rect 551 58 558 60
rect 564 63 571 65
rect 564 61 566 63
rect 568 61 571 63
rect 564 59 571 61
rect 551 50 556 58
rect 531 43 539 50
rect 566 44 571 59
rect 573 62 578 71
rect 595 69 607 71
rect 595 67 602 69
rect 604 67 607 69
rect 595 62 607 67
rect 573 55 581 62
rect 573 53 576 55
rect 578 53 581 55
rect 573 44 581 53
rect 583 55 591 62
rect 583 53 586 55
rect 588 53 591 55
rect 583 48 591 53
rect 583 46 586 48
rect 588 46 591 48
rect 583 44 591 46
rect 593 60 602 62
rect 604 60 607 62
rect 593 44 607 60
rect 609 50 614 71
rect 609 48 616 50
rect 609 46 612 48
rect 614 46 616 48
rect 609 44 616 46
<< alu1 >>
rect 2 288 632 293
rect 2 286 9 288
rect 11 286 58 288
rect 60 286 68 288
rect 70 286 98 288
rect 100 286 151 288
rect 153 286 172 288
rect 174 286 182 288
rect 184 286 212 288
rect 214 286 265 288
rect 267 286 301 288
rect 303 286 311 288
rect 313 286 525 288
rect 527 286 566 288
rect 568 286 619 288
rect 621 286 632 288
rect 2 285 632 286
rect 55 276 67 280
rect 55 274 57 276
rect 59 274 67 276
rect 131 278 155 279
rect 6 271 11 273
rect 6 269 8 271
rect 10 269 11 271
rect 6 267 11 269
rect 6 248 10 267
rect 38 263 42 272
rect 6 246 8 248
rect 6 241 10 246
rect 6 239 8 241
rect 21 262 42 263
rect 21 260 25 262
rect 27 260 39 262
rect 41 260 42 262
rect 21 259 42 260
rect 21 253 35 255
rect 37 253 42 255
rect 21 251 42 253
rect 38 249 42 251
rect 55 254 59 274
rect 131 276 133 278
rect 135 276 155 278
rect 131 275 155 276
rect 79 271 84 272
rect 79 269 80 271
rect 82 269 84 271
rect 79 263 84 269
rect 55 252 60 254
rect 55 250 57 252
rect 59 250 60 252
rect 55 249 60 250
rect 38 245 60 249
rect 38 242 42 245
rect 55 243 57 245
rect 59 243 60 245
rect 70 262 84 263
rect 70 260 74 262
rect 76 260 84 262
rect 70 259 84 260
rect 103 271 116 272
rect 103 269 105 271
rect 107 269 116 271
rect 103 267 116 269
rect 103 266 113 267
rect 111 265 113 266
rect 115 265 116 267
rect 78 254 91 255
rect 78 252 84 254
rect 86 252 91 254
rect 78 251 91 252
rect 55 241 60 243
rect 6 235 19 239
rect 6 234 10 235
rect 87 247 91 251
rect 87 245 88 247
rect 90 245 91 247
rect 87 242 91 245
rect 95 254 100 256
rect 95 252 97 254
rect 99 252 100 254
rect 95 247 100 252
rect 111 258 116 265
rect 151 270 155 275
rect 151 268 152 270
rect 154 268 155 270
rect 95 245 97 247
rect 99 245 100 247
rect 95 240 100 245
rect 95 234 107 240
rect 151 247 155 268
rect 139 245 155 247
rect 139 243 141 245
rect 143 243 155 245
rect 139 242 155 243
rect 169 276 181 280
rect 169 274 171 276
rect 173 274 181 276
rect 245 278 269 279
rect 169 262 173 274
rect 245 276 247 278
rect 249 276 269 278
rect 245 275 269 276
rect 169 260 170 262
rect 172 260 173 262
rect 169 254 173 260
rect 193 271 198 272
rect 193 269 194 271
rect 196 269 198 271
rect 193 263 198 269
rect 169 252 174 254
rect 169 250 171 252
rect 173 250 174 252
rect 169 245 174 250
rect 169 243 171 245
rect 173 243 174 245
rect 184 262 198 263
rect 184 260 188 262
rect 190 260 198 262
rect 184 259 198 260
rect 217 271 230 272
rect 217 269 219 271
rect 221 269 230 271
rect 217 267 230 269
rect 217 266 227 267
rect 225 265 227 266
rect 229 265 230 267
rect 192 254 205 255
rect 192 252 198 254
rect 200 252 205 254
rect 192 251 205 252
rect 169 241 174 243
rect 201 247 205 251
rect 201 245 202 247
rect 204 245 205 247
rect 201 242 205 245
rect 209 254 214 256
rect 209 252 211 254
rect 213 252 214 254
rect 209 247 214 252
rect 225 258 230 265
rect 209 245 211 247
rect 213 245 214 247
rect 209 240 214 245
rect 209 234 221 240
rect 265 255 269 275
rect 287 263 292 272
rect 304 276 316 280
rect 304 274 312 276
rect 314 274 316 276
rect 287 262 301 263
rect 287 260 295 262
rect 297 260 301 262
rect 287 259 301 260
rect 265 253 266 255
rect 268 253 269 255
rect 265 247 269 253
rect 253 245 269 247
rect 253 243 255 245
rect 257 243 269 245
rect 253 242 269 243
rect 280 254 293 255
rect 280 252 285 254
rect 287 252 293 254
rect 280 251 293 252
rect 280 242 284 251
rect 312 270 316 274
rect 312 268 313 270
rect 315 268 316 270
rect 312 254 316 268
rect 311 252 316 254
rect 311 250 312 252
rect 314 250 316 252
rect 378 278 382 280
rect 377 276 382 278
rect 377 274 378 276
rect 380 274 382 276
rect 377 272 382 274
rect 329 270 342 271
rect 329 268 330 270
rect 332 268 342 270
rect 329 267 342 268
rect 336 262 342 267
rect 336 260 337 262
rect 339 260 342 262
rect 336 258 342 260
rect 362 257 366 264
rect 362 256 364 257
rect 354 255 364 256
rect 354 254 366 255
rect 354 252 355 254
rect 357 252 366 254
rect 354 250 366 252
rect 311 245 316 250
rect 311 243 312 245
rect 314 243 316 245
rect 311 241 316 243
rect 322 246 335 247
rect 322 244 332 246
rect 334 244 335 246
rect 322 243 335 244
rect 322 242 327 243
rect 378 262 382 272
rect 378 260 379 262
rect 381 260 382 262
rect 322 240 324 242
rect 326 240 327 242
rect 322 234 327 240
rect 378 239 382 260
rect 369 238 382 239
rect 369 236 378 238
rect 380 236 382 238
rect 369 235 382 236
rect 389 278 393 280
rect 389 276 394 278
rect 389 274 391 276
rect 393 274 394 276
rect 456 278 460 280
rect 389 272 394 274
rect 389 239 393 272
rect 429 270 442 271
rect 405 262 409 264
rect 405 260 406 262
rect 408 260 409 262
rect 405 257 409 260
rect 407 256 409 257
rect 407 255 417 256
rect 405 250 417 255
rect 429 268 437 270
rect 439 268 442 270
rect 429 267 442 268
rect 429 262 435 267
rect 429 260 432 262
rect 434 260 435 262
rect 429 258 435 260
rect 456 276 461 278
rect 456 274 458 276
rect 460 274 461 276
rect 564 278 588 279
rect 456 272 461 274
rect 456 270 460 272
rect 456 268 457 270
rect 459 268 460 270
rect 496 270 509 271
rect 436 243 449 247
rect 444 242 449 243
rect 389 238 402 239
rect 444 240 445 242
rect 447 240 449 242
rect 389 236 391 238
rect 393 236 402 238
rect 389 235 402 236
rect 444 234 449 240
rect 456 239 460 268
rect 472 257 476 264
rect 474 256 476 257
rect 474 255 484 256
rect 472 253 480 255
rect 482 253 484 255
rect 472 250 484 253
rect 496 268 505 270
rect 507 268 509 270
rect 496 267 509 268
rect 496 262 502 267
rect 496 260 499 262
rect 501 260 502 262
rect 496 258 502 260
rect 564 276 584 278
rect 586 276 588 278
rect 564 275 588 276
rect 522 271 527 273
rect 522 269 524 271
rect 526 269 527 271
rect 522 267 527 269
rect 522 254 526 267
rect 522 252 523 254
rect 525 252 526 254
rect 522 248 526 252
rect 554 263 558 272
rect 503 246 516 247
rect 503 244 504 246
rect 506 244 516 246
rect 503 243 516 244
rect 511 242 516 243
rect 456 238 469 239
rect 511 240 512 242
rect 514 240 516 242
rect 456 236 458 238
rect 460 236 469 238
rect 456 235 469 236
rect 511 234 516 240
rect 522 246 524 248
rect 522 241 526 246
rect 522 239 524 241
rect 537 262 558 263
rect 537 260 541 262
rect 543 260 558 262
rect 537 259 558 260
rect 564 270 568 275
rect 564 268 565 270
rect 567 268 568 270
rect 537 253 551 255
rect 553 253 558 255
rect 537 251 558 253
rect 554 242 558 251
rect 564 247 568 268
rect 603 267 616 272
rect 603 265 604 267
rect 606 266 616 267
rect 606 265 608 266
rect 564 245 580 247
rect 564 243 576 245
rect 578 243 580 245
rect 564 242 580 243
rect 603 258 608 265
rect 619 254 624 256
rect 619 252 620 254
rect 622 252 624 254
rect 522 235 535 239
rect 619 240 624 252
rect 522 234 526 235
rect 612 234 624 240
rect 2 228 632 229
rect 2 226 9 228
rect 11 226 58 228
rect 60 226 131 228
rect 133 226 172 228
rect 174 226 245 228
rect 247 226 311 228
rect 313 226 525 228
rect 527 226 586 228
rect 588 226 632 228
rect 2 216 632 226
rect 2 214 9 216
rect 11 214 58 216
rect 60 214 131 216
rect 133 214 172 216
rect 174 214 245 216
rect 247 214 311 216
rect 313 214 525 216
rect 527 214 586 216
rect 588 214 632 216
rect 2 213 632 214
rect 6 207 10 208
rect 6 203 19 207
rect 6 201 8 203
rect 6 196 10 201
rect 6 194 8 196
rect 6 175 10 194
rect 38 197 42 200
rect 55 199 60 201
rect 55 197 57 199
rect 59 197 60 199
rect 95 202 107 208
rect 38 193 60 197
rect 38 191 42 193
rect 21 189 42 191
rect 21 187 35 189
rect 37 187 42 189
rect 55 192 60 193
rect 55 190 57 192
rect 59 190 60 192
rect 55 188 60 190
rect 87 197 91 200
rect 87 195 88 197
rect 90 195 91 197
rect 6 173 11 175
rect 6 171 8 173
rect 10 171 11 173
rect 6 169 11 171
rect 21 182 42 183
rect 21 180 25 182
rect 27 180 39 182
rect 41 180 42 182
rect 21 179 42 180
rect 38 170 42 179
rect 55 168 59 188
rect 87 191 91 195
rect 78 190 91 191
rect 78 188 84 190
rect 86 188 91 190
rect 78 187 91 188
rect 95 197 100 202
rect 95 195 97 197
rect 99 195 100 197
rect 95 190 100 195
rect 95 188 97 190
rect 99 188 100 190
rect 95 186 100 188
rect 70 182 84 183
rect 70 180 74 182
rect 76 180 84 182
rect 70 179 84 180
rect 55 166 57 168
rect 59 166 67 168
rect 55 162 67 166
rect 79 173 84 179
rect 79 171 80 173
rect 82 171 84 173
rect 79 170 84 171
rect 111 177 116 184
rect 139 199 155 200
rect 139 197 141 199
rect 143 197 155 199
rect 139 195 155 197
rect 111 176 113 177
rect 103 175 113 176
rect 115 175 116 177
rect 103 173 116 175
rect 103 171 105 173
rect 107 171 116 173
rect 103 170 116 171
rect 151 174 155 195
rect 151 172 152 174
rect 154 172 155 174
rect 151 167 155 172
rect 131 166 155 167
rect 131 164 133 166
rect 135 164 155 166
rect 131 163 155 164
rect 169 199 174 201
rect 169 197 171 199
rect 173 197 174 199
rect 209 202 221 208
rect 169 192 174 197
rect 169 190 171 192
rect 173 190 174 192
rect 169 188 174 190
rect 201 197 205 200
rect 201 195 202 197
rect 204 195 205 197
rect 169 182 173 188
rect 169 180 170 182
rect 172 180 173 182
rect 169 168 173 180
rect 201 191 205 195
rect 192 190 205 191
rect 192 188 198 190
rect 200 188 205 190
rect 192 187 205 188
rect 209 197 214 202
rect 209 195 211 197
rect 213 195 214 197
rect 209 190 214 195
rect 209 188 211 190
rect 213 188 214 190
rect 209 186 214 188
rect 184 182 198 183
rect 184 180 188 182
rect 190 180 198 182
rect 184 179 198 180
rect 169 166 171 168
rect 173 166 181 168
rect 169 162 181 166
rect 193 173 198 179
rect 193 171 194 173
rect 196 171 198 173
rect 193 170 198 171
rect 225 177 230 184
rect 253 199 269 200
rect 253 197 255 199
rect 257 197 269 199
rect 253 195 269 197
rect 265 189 269 195
rect 265 187 266 189
rect 268 187 269 189
rect 280 191 284 200
rect 322 202 327 208
rect 369 206 382 207
rect 369 204 378 206
rect 380 204 382 206
rect 311 199 316 201
rect 280 190 293 191
rect 280 188 285 190
rect 287 188 293 190
rect 280 187 293 188
rect 225 176 227 177
rect 217 175 227 176
rect 229 175 230 177
rect 217 173 230 175
rect 217 171 219 173
rect 221 171 230 173
rect 217 170 230 171
rect 265 167 269 187
rect 287 182 301 183
rect 287 180 295 182
rect 297 180 301 182
rect 287 179 301 180
rect 311 197 312 199
rect 314 197 316 199
rect 311 192 316 197
rect 322 200 324 202
rect 326 200 327 202
rect 369 203 382 204
rect 322 199 327 200
rect 322 198 335 199
rect 322 196 332 198
rect 334 196 335 198
rect 322 195 335 196
rect 311 190 312 192
rect 314 190 316 192
rect 311 188 316 190
rect 287 170 292 179
rect 312 174 316 188
rect 312 172 313 174
rect 315 172 316 174
rect 312 168 316 172
rect 245 166 269 167
rect 245 164 247 166
rect 249 164 269 166
rect 245 163 269 164
rect 304 166 312 168
rect 314 166 316 168
rect 304 162 316 166
rect 336 182 342 184
rect 336 180 337 182
rect 339 180 342 182
rect 336 175 342 180
rect 329 174 342 175
rect 329 172 330 174
rect 332 172 342 174
rect 354 190 366 192
rect 354 188 355 190
rect 357 188 366 190
rect 354 187 366 188
rect 354 186 364 187
rect 362 185 364 186
rect 362 178 366 185
rect 378 182 382 203
rect 378 180 379 182
rect 381 180 382 182
rect 329 171 342 172
rect 378 170 382 180
rect 377 168 382 170
rect 377 166 378 168
rect 380 166 382 168
rect 377 164 382 166
rect 378 162 382 164
rect 389 206 402 207
rect 389 204 391 206
rect 393 204 402 206
rect 389 203 402 204
rect 389 170 393 203
rect 444 202 449 208
rect 444 200 445 202
rect 447 200 449 202
rect 444 199 449 200
rect 436 195 449 199
rect 456 206 469 207
rect 456 204 458 206
rect 460 204 469 206
rect 456 203 469 204
rect 405 187 417 192
rect 407 186 417 187
rect 407 185 409 186
rect 405 182 409 185
rect 405 180 406 182
rect 408 180 409 182
rect 405 178 409 180
rect 429 182 435 184
rect 429 180 432 182
rect 434 180 435 182
rect 429 175 435 180
rect 429 174 442 175
rect 429 172 437 174
rect 439 172 442 174
rect 429 171 442 172
rect 389 168 394 170
rect 389 166 391 168
rect 393 166 394 168
rect 389 164 394 166
rect 389 162 393 164
rect 456 174 460 203
rect 511 202 516 208
rect 511 200 512 202
rect 514 200 516 202
rect 511 199 516 200
rect 503 198 516 199
rect 503 196 504 198
rect 506 196 516 198
rect 503 195 516 196
rect 522 207 526 208
rect 522 203 535 207
rect 522 201 524 203
rect 522 196 526 201
rect 522 194 524 196
rect 472 189 484 192
rect 472 187 480 189
rect 482 187 484 189
rect 474 186 484 187
rect 474 185 476 186
rect 456 172 457 174
rect 459 172 460 174
rect 472 178 476 185
rect 456 170 460 172
rect 496 182 502 184
rect 496 180 499 182
rect 501 180 502 182
rect 496 175 502 180
rect 496 174 509 175
rect 496 172 505 174
rect 507 172 509 174
rect 496 171 509 172
rect 456 168 461 170
rect 456 166 458 168
rect 460 166 461 168
rect 456 164 461 166
rect 456 162 460 164
rect 522 190 526 194
rect 522 188 523 190
rect 525 188 526 190
rect 522 175 526 188
rect 554 191 558 200
rect 537 189 558 191
rect 537 187 551 189
rect 553 187 558 189
rect 564 199 580 200
rect 564 197 576 199
rect 578 197 580 199
rect 564 195 580 197
rect 522 173 527 175
rect 522 171 524 173
rect 526 171 527 173
rect 522 169 527 171
rect 537 182 558 183
rect 537 180 541 182
rect 543 180 558 182
rect 537 179 558 180
rect 554 170 558 179
rect 564 174 568 195
rect 612 202 624 208
rect 564 172 565 174
rect 567 172 568 174
rect 564 167 568 172
rect 603 177 608 184
rect 619 190 624 202
rect 619 188 620 190
rect 622 188 624 190
rect 619 186 624 188
rect 603 175 604 177
rect 606 176 608 177
rect 606 175 616 176
rect 603 170 616 175
rect 564 166 588 167
rect 564 164 584 166
rect 586 164 588 166
rect 564 163 588 164
rect 2 156 632 157
rect 2 154 9 156
rect 11 154 58 156
rect 60 154 68 156
rect 70 154 98 156
rect 100 154 151 156
rect 153 154 172 156
rect 174 154 182 156
rect 184 154 212 156
rect 214 154 265 156
rect 267 154 301 156
rect 303 154 311 156
rect 313 154 525 156
rect 527 154 566 156
rect 568 154 619 156
rect 621 154 632 156
rect 2 144 632 154
rect 2 142 9 144
rect 11 142 58 144
rect 60 142 68 144
rect 70 142 98 144
rect 100 142 151 144
rect 153 142 172 144
rect 174 142 182 144
rect 184 142 212 144
rect 214 142 265 144
rect 267 142 301 144
rect 303 142 311 144
rect 313 142 525 144
rect 527 142 566 144
rect 568 142 619 144
rect 621 142 632 144
rect 2 141 632 142
rect 55 132 67 136
rect 55 130 57 132
rect 59 130 67 132
rect 131 134 155 135
rect 6 127 11 129
rect 6 125 8 127
rect 10 125 11 127
rect 6 123 11 125
rect 6 104 10 123
rect 38 119 42 128
rect 6 102 8 104
rect 6 97 10 102
rect 6 95 8 97
rect 21 118 42 119
rect 21 116 25 118
rect 27 116 39 118
rect 41 116 42 118
rect 21 115 42 116
rect 21 109 35 111
rect 37 109 42 111
rect 21 107 42 109
rect 38 105 42 107
rect 55 110 59 130
rect 131 132 133 134
rect 135 132 155 134
rect 131 131 155 132
rect 79 127 84 128
rect 79 125 80 127
rect 82 125 84 127
rect 79 119 84 125
rect 55 108 60 110
rect 55 106 57 108
rect 59 106 60 108
rect 55 105 60 106
rect 38 101 60 105
rect 38 98 42 101
rect 55 99 57 101
rect 59 99 60 101
rect 70 118 84 119
rect 70 116 74 118
rect 76 116 84 118
rect 70 115 84 116
rect 103 127 116 128
rect 103 125 105 127
rect 107 125 116 127
rect 103 123 116 125
rect 103 122 113 123
rect 111 121 113 122
rect 115 121 116 123
rect 78 110 91 111
rect 78 108 84 110
rect 86 108 91 110
rect 78 107 91 108
rect 55 97 60 99
rect 6 91 19 95
rect 6 90 10 91
rect 87 103 91 107
rect 87 101 88 103
rect 90 101 91 103
rect 87 98 91 101
rect 95 110 100 112
rect 95 108 97 110
rect 99 108 100 110
rect 95 103 100 108
rect 111 114 116 121
rect 151 126 155 131
rect 151 124 152 126
rect 154 124 155 126
rect 95 101 97 103
rect 99 101 100 103
rect 95 96 100 101
rect 95 90 107 96
rect 151 103 155 124
rect 139 101 155 103
rect 139 99 141 101
rect 143 99 155 101
rect 139 98 155 99
rect 169 132 181 136
rect 169 130 171 132
rect 173 130 181 132
rect 245 134 269 135
rect 169 118 173 130
rect 245 132 247 134
rect 249 132 269 134
rect 245 131 269 132
rect 169 116 170 118
rect 172 116 173 118
rect 169 110 173 116
rect 193 127 198 128
rect 193 125 194 127
rect 196 125 198 127
rect 193 119 198 125
rect 169 108 174 110
rect 169 106 171 108
rect 173 106 174 108
rect 169 101 174 106
rect 169 99 171 101
rect 173 99 174 101
rect 184 118 198 119
rect 184 116 188 118
rect 190 116 198 118
rect 184 115 198 116
rect 217 127 230 128
rect 217 125 219 127
rect 221 125 230 127
rect 217 123 230 125
rect 217 122 227 123
rect 225 121 227 122
rect 229 121 230 123
rect 192 110 205 111
rect 192 108 198 110
rect 200 108 205 110
rect 192 107 205 108
rect 169 97 174 99
rect 201 103 205 107
rect 201 101 202 103
rect 204 101 205 103
rect 201 98 205 101
rect 209 110 214 112
rect 209 108 211 110
rect 213 108 214 110
rect 209 103 214 108
rect 225 114 230 121
rect 209 101 211 103
rect 213 101 214 103
rect 209 96 214 101
rect 209 90 221 96
rect 265 111 269 131
rect 287 119 292 128
rect 304 132 316 136
rect 304 130 312 132
rect 314 130 316 132
rect 287 118 301 119
rect 287 116 295 118
rect 297 116 301 118
rect 287 115 301 116
rect 265 109 266 111
rect 268 109 269 111
rect 265 103 269 109
rect 253 101 269 103
rect 253 99 255 101
rect 257 99 269 101
rect 253 98 269 99
rect 280 110 293 111
rect 280 108 285 110
rect 287 108 293 110
rect 280 107 293 108
rect 280 98 284 107
rect 312 126 316 130
rect 312 124 313 126
rect 315 124 316 126
rect 312 110 316 124
rect 311 108 316 110
rect 311 106 312 108
rect 314 106 316 108
rect 378 134 382 136
rect 377 132 382 134
rect 377 130 378 132
rect 380 130 382 132
rect 377 128 382 130
rect 329 126 342 127
rect 329 124 330 126
rect 332 124 342 126
rect 329 123 342 124
rect 336 118 342 123
rect 336 116 337 118
rect 339 116 342 118
rect 336 114 342 116
rect 362 113 366 120
rect 362 112 364 113
rect 354 111 364 112
rect 354 110 366 111
rect 354 108 355 110
rect 357 108 366 110
rect 354 106 366 108
rect 311 101 316 106
rect 311 99 312 101
rect 314 99 316 101
rect 311 97 316 99
rect 322 102 335 103
rect 322 100 332 102
rect 334 100 335 102
rect 322 99 335 100
rect 322 98 327 99
rect 378 118 382 128
rect 378 116 379 118
rect 381 116 382 118
rect 322 96 324 98
rect 326 96 327 98
rect 322 90 327 96
rect 378 95 382 116
rect 369 94 382 95
rect 369 92 378 94
rect 380 92 382 94
rect 369 91 382 92
rect 389 134 393 136
rect 389 132 394 134
rect 389 130 391 132
rect 393 130 394 132
rect 456 134 460 136
rect 389 128 394 130
rect 389 95 393 128
rect 429 126 442 127
rect 405 118 409 120
rect 405 116 406 118
rect 408 116 409 118
rect 405 113 409 116
rect 407 112 409 113
rect 407 111 417 112
rect 405 106 417 111
rect 429 124 437 126
rect 439 124 442 126
rect 429 123 442 124
rect 429 118 435 123
rect 429 116 432 118
rect 434 116 435 118
rect 429 114 435 116
rect 456 132 461 134
rect 456 130 458 132
rect 460 130 461 132
rect 564 134 588 135
rect 456 128 461 130
rect 456 126 460 128
rect 456 124 457 126
rect 459 124 460 126
rect 496 126 509 127
rect 436 99 449 103
rect 444 98 449 99
rect 389 94 402 95
rect 444 96 445 98
rect 447 96 449 98
rect 389 92 391 94
rect 393 92 402 94
rect 389 91 402 92
rect 444 90 449 96
rect 456 95 460 124
rect 472 113 476 120
rect 474 112 476 113
rect 474 111 484 112
rect 472 109 480 111
rect 482 109 484 111
rect 472 106 484 109
rect 496 124 505 126
rect 507 124 509 126
rect 496 123 509 124
rect 496 118 502 123
rect 496 116 499 118
rect 501 116 502 118
rect 496 114 502 116
rect 564 132 584 134
rect 586 132 588 134
rect 564 131 588 132
rect 522 127 527 129
rect 522 125 524 127
rect 526 125 527 127
rect 522 123 527 125
rect 522 110 526 123
rect 522 108 523 110
rect 525 108 526 110
rect 522 104 526 108
rect 554 119 558 128
rect 503 102 516 103
rect 503 100 504 102
rect 506 100 516 102
rect 503 99 516 100
rect 511 98 516 99
rect 456 94 469 95
rect 511 96 512 98
rect 514 96 516 98
rect 456 92 458 94
rect 460 92 469 94
rect 456 91 469 92
rect 511 90 516 96
rect 522 102 524 104
rect 522 97 526 102
rect 522 95 524 97
rect 537 118 558 119
rect 537 116 541 118
rect 543 116 558 118
rect 537 115 558 116
rect 564 126 568 131
rect 564 124 565 126
rect 567 124 568 126
rect 537 109 551 111
rect 553 109 558 111
rect 537 107 558 109
rect 554 98 558 107
rect 564 103 568 124
rect 603 123 616 128
rect 603 121 604 123
rect 606 122 616 123
rect 606 121 608 122
rect 564 101 580 103
rect 564 99 576 101
rect 578 99 580 101
rect 564 98 580 99
rect 603 114 608 121
rect 619 110 624 112
rect 619 108 620 110
rect 622 108 624 110
rect 522 91 535 95
rect 619 96 624 108
rect 522 90 526 91
rect 612 90 624 96
rect 2 84 632 85
rect 2 82 9 84
rect 11 82 58 84
rect 60 82 131 84
rect 133 82 172 84
rect 174 82 245 84
rect 247 82 311 84
rect 313 82 525 84
rect 527 82 586 84
rect 588 82 632 84
rect 2 72 632 82
rect 2 70 9 72
rect 11 70 58 72
rect 60 70 131 72
rect 133 70 172 72
rect 174 70 245 72
rect 247 70 311 72
rect 313 70 525 72
rect 527 70 586 72
rect 588 70 632 72
rect 2 69 632 70
rect 6 63 10 64
rect 6 59 19 63
rect 6 57 8 59
rect 6 52 10 57
rect 6 50 8 52
rect 6 31 10 50
rect 38 53 42 56
rect 55 55 60 57
rect 55 53 57 55
rect 59 53 60 55
rect 95 58 107 64
rect 38 49 60 53
rect 38 47 42 49
rect 21 45 42 47
rect 21 43 35 45
rect 37 43 42 45
rect 55 48 60 49
rect 55 46 57 48
rect 59 46 60 48
rect 55 44 60 46
rect 87 53 91 56
rect 87 51 88 53
rect 90 51 91 53
rect 6 29 11 31
rect 6 27 8 29
rect 10 27 11 29
rect 6 25 11 27
rect 21 38 42 39
rect 21 36 25 38
rect 27 36 39 38
rect 41 36 42 38
rect 21 35 42 36
rect 38 26 42 35
rect 55 24 59 44
rect 87 47 91 51
rect 78 46 91 47
rect 78 44 84 46
rect 86 44 91 46
rect 78 43 91 44
rect 95 53 100 58
rect 95 51 97 53
rect 99 51 100 53
rect 95 46 100 51
rect 95 44 97 46
rect 99 44 100 46
rect 95 42 100 44
rect 70 38 84 39
rect 70 36 74 38
rect 76 36 84 38
rect 70 35 84 36
rect 55 22 57 24
rect 59 22 67 24
rect 55 18 67 22
rect 79 29 84 35
rect 79 27 80 29
rect 82 27 84 29
rect 79 26 84 27
rect 111 33 116 40
rect 139 55 155 56
rect 139 53 141 55
rect 143 53 155 55
rect 139 51 155 53
rect 111 32 113 33
rect 103 31 113 32
rect 115 31 116 33
rect 103 29 116 31
rect 103 27 105 29
rect 107 27 116 29
rect 103 26 116 27
rect 151 30 155 51
rect 151 28 152 30
rect 154 28 155 30
rect 151 23 155 28
rect 131 22 155 23
rect 131 20 133 22
rect 135 20 155 22
rect 131 19 155 20
rect 169 55 174 57
rect 169 53 171 55
rect 173 53 174 55
rect 209 58 221 64
rect 169 48 174 53
rect 169 46 171 48
rect 173 46 174 48
rect 169 44 174 46
rect 201 53 205 56
rect 201 51 202 53
rect 204 51 205 53
rect 169 38 173 44
rect 169 36 170 38
rect 172 36 173 38
rect 169 24 173 36
rect 201 47 205 51
rect 192 46 205 47
rect 192 44 198 46
rect 200 44 205 46
rect 192 43 205 44
rect 209 53 214 58
rect 209 51 211 53
rect 213 51 214 53
rect 209 46 214 51
rect 209 44 211 46
rect 213 44 214 46
rect 209 42 214 44
rect 184 38 198 39
rect 184 36 188 38
rect 190 36 198 38
rect 184 35 198 36
rect 169 22 171 24
rect 173 22 181 24
rect 169 18 181 22
rect 193 29 198 35
rect 193 27 194 29
rect 196 27 198 29
rect 193 26 198 27
rect 225 33 230 40
rect 253 55 269 56
rect 253 53 255 55
rect 257 53 269 55
rect 253 51 269 53
rect 265 45 269 51
rect 265 43 266 45
rect 268 43 269 45
rect 280 47 284 56
rect 322 58 327 64
rect 369 62 382 63
rect 369 60 378 62
rect 380 60 382 62
rect 311 55 316 57
rect 280 46 293 47
rect 280 44 285 46
rect 287 44 293 46
rect 280 43 293 44
rect 225 32 227 33
rect 217 31 227 32
rect 229 31 230 33
rect 217 29 230 31
rect 217 27 219 29
rect 221 27 230 29
rect 217 26 230 27
rect 265 23 269 43
rect 287 38 301 39
rect 287 36 295 38
rect 297 36 301 38
rect 287 35 301 36
rect 311 53 312 55
rect 314 53 316 55
rect 311 48 316 53
rect 322 56 324 58
rect 326 56 327 58
rect 369 59 382 60
rect 322 55 327 56
rect 322 54 335 55
rect 322 52 332 54
rect 334 52 335 54
rect 322 51 335 52
rect 311 46 312 48
rect 314 46 316 48
rect 311 44 316 46
rect 287 26 292 35
rect 312 30 316 44
rect 312 28 313 30
rect 315 28 316 30
rect 312 24 316 28
rect 245 22 269 23
rect 245 20 247 22
rect 249 20 269 22
rect 245 19 269 20
rect 304 22 312 24
rect 314 22 316 24
rect 304 18 316 22
rect 336 38 342 40
rect 336 36 337 38
rect 339 36 342 38
rect 336 31 342 36
rect 329 30 342 31
rect 329 28 330 30
rect 332 28 342 30
rect 354 46 366 48
rect 354 44 355 46
rect 357 44 366 46
rect 354 43 366 44
rect 354 42 364 43
rect 362 41 364 42
rect 362 34 366 41
rect 378 38 382 59
rect 378 36 379 38
rect 381 36 382 38
rect 329 27 342 28
rect 378 26 382 36
rect 377 24 382 26
rect 377 22 378 24
rect 380 22 382 24
rect 377 20 382 22
rect 378 18 382 20
rect 389 62 402 63
rect 389 60 391 62
rect 393 60 402 62
rect 389 59 402 60
rect 389 26 393 59
rect 444 58 449 64
rect 444 56 445 58
rect 447 56 449 58
rect 444 55 449 56
rect 436 51 449 55
rect 456 62 469 63
rect 456 60 458 62
rect 460 60 469 62
rect 456 59 469 60
rect 405 43 417 48
rect 407 42 417 43
rect 407 41 409 42
rect 405 38 409 41
rect 405 36 406 38
rect 408 36 409 38
rect 405 34 409 36
rect 429 38 435 40
rect 429 36 432 38
rect 434 36 435 38
rect 429 31 435 36
rect 429 30 442 31
rect 429 28 437 30
rect 439 28 442 30
rect 429 27 442 28
rect 389 24 394 26
rect 389 22 391 24
rect 393 22 394 24
rect 389 20 394 22
rect 389 18 393 20
rect 456 30 460 59
rect 511 58 516 64
rect 511 56 512 58
rect 514 56 516 58
rect 511 55 516 56
rect 503 54 516 55
rect 503 52 504 54
rect 506 52 516 54
rect 503 51 516 52
rect 522 63 526 64
rect 522 59 535 63
rect 522 57 524 59
rect 522 52 526 57
rect 522 50 524 52
rect 472 45 484 48
rect 472 43 480 45
rect 482 43 484 45
rect 474 42 484 43
rect 474 41 476 42
rect 456 28 457 30
rect 459 28 460 30
rect 472 34 476 41
rect 456 26 460 28
rect 496 38 502 40
rect 496 36 499 38
rect 501 36 502 38
rect 496 31 502 36
rect 496 30 509 31
rect 496 28 505 30
rect 507 28 509 30
rect 496 27 509 28
rect 456 24 461 26
rect 456 22 458 24
rect 460 22 461 24
rect 456 20 461 22
rect 456 18 460 20
rect 522 46 526 50
rect 522 44 523 46
rect 525 44 526 46
rect 522 31 526 44
rect 554 47 558 56
rect 537 45 558 47
rect 537 43 551 45
rect 553 43 558 45
rect 564 55 580 56
rect 564 53 576 55
rect 578 53 580 55
rect 564 51 580 53
rect 522 29 527 31
rect 522 27 524 29
rect 526 27 527 29
rect 522 25 527 27
rect 537 38 558 39
rect 537 36 541 38
rect 543 36 558 38
rect 537 35 558 36
rect 554 26 558 35
rect 564 30 568 51
rect 612 58 624 64
rect 564 28 565 30
rect 567 28 568 30
rect 564 23 568 28
rect 603 33 608 40
rect 619 46 624 58
rect 619 44 620 46
rect 622 44 624 46
rect 619 42 624 44
rect 603 31 604 33
rect 606 32 608 33
rect 606 31 616 32
rect 603 26 616 31
rect 564 22 588 23
rect 564 20 584 22
rect 586 20 588 22
rect 564 19 588 20
rect 2 12 632 13
rect 2 10 9 12
rect 11 10 58 12
rect 60 10 68 12
rect 70 10 98 12
rect 100 10 151 12
rect 153 10 172 12
rect 174 10 182 12
rect 184 10 212 12
rect 214 10 265 12
rect 267 10 301 12
rect 303 10 311 12
rect 313 10 525 12
rect 527 10 566 12
rect 568 10 619 12
rect 621 10 632 12
rect 2 5 632 10
<< alu2 >>
rect 79 271 111 272
rect 79 269 80 271
rect 82 269 105 271
rect 107 269 111 271
rect 79 267 111 269
rect 151 271 225 272
rect 151 270 194 271
rect 151 268 152 270
rect 154 269 194 270
rect 196 269 219 271
rect 221 269 225 271
rect 154 268 225 269
rect 151 267 225 268
rect 312 270 333 271
rect 312 268 313 270
rect 315 268 330 270
rect 332 268 333 270
rect 312 267 333 268
rect 436 270 460 271
rect 436 268 437 270
rect 439 268 457 270
rect 459 268 460 270
rect 436 267 460 268
rect 504 270 568 271
rect 504 268 505 270
rect 507 268 565 270
rect 567 268 568 270
rect 504 267 568 268
rect 38 262 173 263
rect 38 260 39 262
rect 41 260 170 262
rect 172 260 173 262
rect 38 259 173 260
rect 378 262 409 263
rect 378 260 379 262
rect 381 260 406 262
rect 408 260 409 262
rect 378 259 409 260
rect 265 255 359 256
rect 265 253 266 255
rect 268 254 359 255
rect 268 253 355 254
rect 265 252 355 253
rect 357 252 359 254
rect 265 251 359 252
rect 479 255 526 256
rect 479 253 480 255
rect 482 254 526 255
rect 482 253 523 254
rect 479 252 523 253
rect 525 252 526 254
rect 479 251 526 252
rect 87 247 100 248
rect 87 245 88 247
rect 90 245 97 247
rect 99 245 100 247
rect 87 244 100 245
rect 201 247 214 248
rect 201 245 202 247
rect 204 245 211 247
rect 213 245 214 247
rect 201 244 214 245
rect 331 246 508 247
rect 331 244 332 246
rect 334 244 504 246
rect 506 244 508 246
rect 331 243 508 244
rect 331 198 508 199
rect 87 197 100 198
rect 87 195 88 197
rect 90 195 97 197
rect 99 195 100 197
rect 87 194 100 195
rect 201 197 214 198
rect 201 195 202 197
rect 204 195 211 197
rect 213 195 214 197
rect 331 196 332 198
rect 334 196 504 198
rect 506 196 508 198
rect 331 195 508 196
rect 201 194 214 195
rect 265 190 359 191
rect 265 189 355 190
rect 265 187 266 189
rect 268 188 355 189
rect 357 188 359 190
rect 268 187 359 188
rect 265 186 359 187
rect 479 190 526 191
rect 479 189 523 190
rect 479 187 480 189
rect 482 188 523 189
rect 525 188 526 190
rect 482 187 526 188
rect 479 186 526 187
rect 38 182 173 183
rect 38 180 39 182
rect 41 180 170 182
rect 172 180 173 182
rect 38 179 173 180
rect 378 182 409 183
rect 378 180 379 182
rect 381 180 406 182
rect 408 180 409 182
rect 378 179 409 180
rect 79 173 111 175
rect 79 171 80 173
rect 82 171 105 173
rect 107 171 111 173
rect 79 170 111 171
rect 151 174 225 175
rect 151 172 152 174
rect 154 173 225 174
rect 154 172 194 173
rect 151 171 194 172
rect 196 171 219 173
rect 221 171 225 173
rect 312 174 333 175
rect 312 172 313 174
rect 315 172 330 174
rect 332 172 333 174
rect 312 171 333 172
rect 436 174 460 175
rect 436 172 437 174
rect 439 172 457 174
rect 459 172 460 174
rect 436 171 460 172
rect 504 174 568 175
rect 504 172 505 174
rect 507 172 565 174
rect 567 172 568 174
rect 504 171 568 172
rect 151 170 225 171
rect 79 127 111 128
rect 79 125 80 127
rect 82 125 105 127
rect 107 125 111 127
rect 79 123 111 125
rect 151 127 225 128
rect 151 126 194 127
rect 151 124 152 126
rect 154 125 194 126
rect 196 125 219 127
rect 221 125 225 127
rect 154 124 225 125
rect 151 123 225 124
rect 312 126 333 127
rect 312 124 313 126
rect 315 124 330 126
rect 332 124 333 126
rect 312 123 333 124
rect 436 126 460 127
rect 436 124 437 126
rect 439 124 457 126
rect 459 124 460 126
rect 436 123 460 124
rect 504 126 568 127
rect 504 124 505 126
rect 507 124 565 126
rect 567 124 568 126
rect 504 123 568 124
rect 38 118 173 119
rect 38 116 39 118
rect 41 116 170 118
rect 172 116 173 118
rect 38 115 173 116
rect 378 118 409 119
rect 378 116 379 118
rect 381 116 406 118
rect 408 116 409 118
rect 378 115 409 116
rect 265 111 359 112
rect 265 109 266 111
rect 268 110 359 111
rect 268 109 355 110
rect 265 108 355 109
rect 357 108 359 110
rect 265 107 359 108
rect 479 111 526 112
rect 479 109 480 111
rect 482 110 526 111
rect 482 109 523 110
rect 479 108 523 109
rect 525 108 526 110
rect 479 107 526 108
rect 87 103 100 104
rect 87 101 88 103
rect 90 101 97 103
rect 99 101 100 103
rect 87 100 100 101
rect 201 103 214 104
rect 201 101 202 103
rect 204 101 211 103
rect 213 101 214 103
rect 201 100 214 101
rect 331 102 508 103
rect 331 100 332 102
rect 334 100 504 102
rect 506 100 508 102
rect 331 99 508 100
rect 331 54 508 55
rect 87 53 100 54
rect 87 51 88 53
rect 90 51 97 53
rect 99 51 100 53
rect 87 50 100 51
rect 201 53 214 54
rect 201 51 202 53
rect 204 51 211 53
rect 213 51 214 53
rect 331 52 332 54
rect 334 52 504 54
rect 506 52 508 54
rect 331 51 508 52
rect 201 50 214 51
rect 265 46 359 47
rect 265 45 355 46
rect 265 43 266 45
rect 268 44 355 45
rect 357 44 359 46
rect 268 43 359 44
rect 265 42 359 43
rect 479 46 526 47
rect 479 45 523 46
rect 479 43 480 45
rect 482 44 523 45
rect 525 44 526 46
rect 482 43 526 44
rect 479 42 526 43
rect 38 38 173 39
rect 38 36 39 38
rect 41 36 170 38
rect 172 36 173 38
rect 38 35 173 36
rect 378 38 409 39
rect 378 36 379 38
rect 381 36 406 38
rect 408 36 409 38
rect 378 35 409 36
rect 79 29 111 31
rect 79 27 80 29
rect 82 27 105 29
rect 107 27 111 29
rect 79 26 111 27
rect 151 30 225 31
rect 151 28 152 30
rect 154 29 225 30
rect 154 28 194 29
rect 151 27 194 28
rect 196 27 219 29
rect 221 27 225 29
rect 312 30 333 31
rect 312 28 313 30
rect 315 28 330 30
rect 332 28 333 30
rect 312 27 333 28
rect 436 30 460 31
rect 436 28 437 30
rect 439 28 457 30
rect 459 28 460 30
rect 436 27 460 28
rect 504 30 568 31
rect 504 28 505 30
rect 507 28 565 30
rect 567 28 568 30
rect 504 27 568 28
rect 151 26 225 27
<< ptie >>
rect 7 288 13 290
rect 7 286 9 288
rect 11 286 13 288
rect 56 288 62 290
rect 56 286 58 288
rect 60 286 62 288
rect 7 284 13 286
rect 56 284 62 286
rect 96 288 102 290
rect 96 286 98 288
rect 100 286 102 288
rect 96 284 102 286
rect 170 288 176 290
rect 170 286 172 288
rect 174 286 176 288
rect 170 284 176 286
rect 210 288 216 290
rect 210 286 212 288
rect 214 286 216 288
rect 210 284 216 286
rect 309 288 315 290
rect 309 286 311 288
rect 313 286 315 288
rect 309 284 315 286
rect 523 288 529 290
rect 523 286 525 288
rect 527 286 529 288
rect 523 284 529 286
rect 617 288 623 290
rect 617 286 619 288
rect 621 286 623 288
rect 617 284 623 286
rect 7 156 13 158
rect 56 156 62 158
rect 7 154 9 156
rect 11 154 13 156
rect 7 152 13 154
rect 56 154 58 156
rect 60 154 62 156
rect 56 152 62 154
rect 96 156 102 158
rect 96 154 98 156
rect 100 154 102 156
rect 96 152 102 154
rect 170 156 176 158
rect 170 154 172 156
rect 174 154 176 156
rect 170 152 176 154
rect 210 156 216 158
rect 210 154 212 156
rect 214 154 216 156
rect 210 152 216 154
rect 309 156 315 158
rect 309 154 311 156
rect 313 154 315 156
rect 309 152 315 154
rect 523 156 529 158
rect 523 154 525 156
rect 527 154 529 156
rect 523 152 529 154
rect 617 156 623 158
rect 617 154 619 156
rect 621 154 623 156
rect 617 152 623 154
rect 7 144 13 146
rect 7 142 9 144
rect 11 142 13 144
rect 56 144 62 146
rect 56 142 58 144
rect 60 142 62 144
rect 7 140 13 142
rect 56 140 62 142
rect 96 144 102 146
rect 96 142 98 144
rect 100 142 102 144
rect 96 140 102 142
rect 170 144 176 146
rect 170 142 172 144
rect 174 142 176 144
rect 170 140 176 142
rect 210 144 216 146
rect 210 142 212 144
rect 214 142 216 144
rect 210 140 216 142
rect 309 144 315 146
rect 309 142 311 144
rect 313 142 315 144
rect 309 140 315 142
rect 523 144 529 146
rect 523 142 525 144
rect 527 142 529 144
rect 523 140 529 142
rect 617 144 623 146
rect 617 142 619 144
rect 621 142 623 144
rect 617 140 623 142
rect 7 12 13 14
rect 56 12 62 14
rect 7 10 9 12
rect 11 10 13 12
rect 7 8 13 10
rect 56 10 58 12
rect 60 10 62 12
rect 56 8 62 10
rect 96 12 102 14
rect 96 10 98 12
rect 100 10 102 12
rect 96 8 102 10
rect 170 12 176 14
rect 170 10 172 12
rect 174 10 176 12
rect 170 8 176 10
rect 210 12 216 14
rect 210 10 212 12
rect 214 10 216 12
rect 210 8 216 10
rect 309 12 315 14
rect 309 10 311 12
rect 313 10 315 12
rect 309 8 315 10
rect 523 12 529 14
rect 523 10 525 12
rect 527 10 529 12
rect 523 8 529 10
rect 617 12 623 14
rect 617 10 619 12
rect 621 10 623 12
rect 617 8 623 10
<< ntie >>
rect 7 228 13 230
rect 7 226 9 228
rect 11 226 13 228
rect 56 228 62 230
rect 7 224 13 226
rect 56 226 58 228
rect 60 226 62 228
rect 129 228 135 230
rect 56 224 62 226
rect 129 226 131 228
rect 133 226 135 228
rect 170 228 176 230
rect 129 224 135 226
rect 170 226 172 228
rect 174 226 176 228
rect 243 228 249 230
rect 170 224 176 226
rect 243 226 245 228
rect 247 226 249 228
rect 309 228 315 230
rect 243 224 249 226
rect 309 226 311 228
rect 313 226 315 228
rect 523 228 529 230
rect 309 224 315 226
rect 523 226 525 228
rect 527 226 529 228
rect 584 228 590 230
rect 523 224 529 226
rect 584 226 586 228
rect 588 226 590 228
rect 584 224 590 226
rect 7 216 13 218
rect 7 214 9 216
rect 11 214 13 216
rect 56 216 62 218
rect 7 212 13 214
rect 56 214 58 216
rect 60 214 62 216
rect 129 216 135 218
rect 56 212 62 214
rect 129 214 131 216
rect 133 214 135 216
rect 170 216 176 218
rect 129 212 135 214
rect 170 214 172 216
rect 174 214 176 216
rect 243 216 249 218
rect 170 212 176 214
rect 243 214 245 216
rect 247 214 249 216
rect 309 216 315 218
rect 243 212 249 214
rect 309 214 311 216
rect 313 214 315 216
rect 523 216 529 218
rect 309 212 315 214
rect 523 214 525 216
rect 527 214 529 216
rect 584 216 590 218
rect 523 212 529 214
rect 584 214 586 216
rect 588 214 590 216
rect 584 212 590 214
rect 7 84 13 86
rect 7 82 9 84
rect 11 82 13 84
rect 56 84 62 86
rect 7 80 13 82
rect 56 82 58 84
rect 60 82 62 84
rect 129 84 135 86
rect 56 80 62 82
rect 129 82 131 84
rect 133 82 135 84
rect 170 84 176 86
rect 129 80 135 82
rect 170 82 172 84
rect 174 82 176 84
rect 243 84 249 86
rect 170 80 176 82
rect 243 82 245 84
rect 247 82 249 84
rect 309 84 315 86
rect 243 80 249 82
rect 309 82 311 84
rect 313 82 315 84
rect 523 84 529 86
rect 309 80 315 82
rect 523 82 525 84
rect 527 82 529 84
rect 584 84 590 86
rect 523 80 529 82
rect 584 82 586 84
rect 588 82 590 84
rect 584 80 590 82
rect 7 72 13 74
rect 7 70 9 72
rect 11 70 13 72
rect 56 72 62 74
rect 7 68 13 70
rect 56 70 58 72
rect 60 70 62 72
rect 129 72 135 74
rect 56 68 62 70
rect 129 70 131 72
rect 133 70 135 72
rect 170 72 176 74
rect 129 68 135 70
rect 170 70 172 72
rect 174 70 176 72
rect 243 72 249 74
rect 170 68 176 70
rect 243 70 245 72
rect 247 70 249 72
rect 309 72 315 74
rect 243 68 249 70
rect 309 70 311 72
rect 313 70 315 72
rect 523 72 529 74
rect 309 68 315 70
rect 523 70 525 72
rect 527 70 529 72
rect 584 72 590 74
rect 523 68 529 70
rect 584 70 586 72
rect 588 70 590 72
rect 584 68 590 70
<< nmos >>
rect 13 267 15 276
rect 23 267 25 273
rect 33 267 35 273
rect 62 269 64 278
rect 75 269 77 280
rect 82 269 84 280
rect 102 267 104 276
rect 118 272 120 281
rect 128 272 130 281
rect 138 272 140 284
rect 145 272 147 284
rect 176 269 178 278
rect 189 269 191 280
rect 196 269 198 280
rect 216 267 218 276
rect 232 272 234 281
rect 242 272 244 281
rect 252 272 254 284
rect 259 272 261 284
rect 287 269 289 280
rect 294 269 296 280
rect 307 269 309 278
rect 329 273 331 279
rect 339 273 341 281
rect 346 273 348 281
rect 356 273 358 281
rect 363 273 365 281
rect 373 272 375 281
rect 396 272 398 281
rect 406 273 408 281
rect 413 273 415 281
rect 423 273 425 281
rect 430 273 432 281
rect 440 273 442 279
rect 463 272 465 281
rect 473 273 475 281
rect 480 273 482 281
rect 490 273 492 281
rect 497 273 499 281
rect 507 273 509 279
rect 529 267 531 276
rect 539 267 541 273
rect 549 267 551 273
rect 572 272 574 284
rect 579 272 581 284
rect 589 272 591 281
rect 599 272 601 281
rect 615 267 617 276
rect 13 166 15 175
rect 23 169 25 175
rect 33 169 35 175
rect 62 164 64 173
rect 75 162 77 173
rect 82 162 84 173
rect 102 166 104 175
rect 118 161 120 170
rect 128 161 130 170
rect 138 158 140 170
rect 145 158 147 170
rect 176 164 178 173
rect 189 162 191 173
rect 196 162 198 173
rect 216 166 218 175
rect 232 161 234 170
rect 242 161 244 170
rect 252 158 254 170
rect 259 158 261 170
rect 287 162 289 173
rect 294 162 296 173
rect 307 164 309 173
rect 329 163 331 169
rect 339 161 341 169
rect 346 161 348 169
rect 356 161 358 169
rect 363 161 365 169
rect 373 161 375 170
rect 396 161 398 170
rect 406 161 408 169
rect 413 161 415 169
rect 423 161 425 169
rect 430 161 432 169
rect 440 163 442 169
rect 463 161 465 170
rect 473 161 475 169
rect 480 161 482 169
rect 490 161 492 169
rect 497 161 499 169
rect 507 163 509 169
rect 529 166 531 175
rect 539 169 541 175
rect 549 169 551 175
rect 572 158 574 170
rect 579 158 581 170
rect 589 161 591 170
rect 599 161 601 170
rect 615 166 617 175
rect 13 123 15 132
rect 23 123 25 129
rect 33 123 35 129
rect 62 125 64 134
rect 75 125 77 136
rect 82 125 84 136
rect 102 123 104 132
rect 118 128 120 137
rect 128 128 130 137
rect 138 128 140 140
rect 145 128 147 140
rect 176 125 178 134
rect 189 125 191 136
rect 196 125 198 136
rect 216 123 218 132
rect 232 128 234 137
rect 242 128 244 137
rect 252 128 254 140
rect 259 128 261 140
rect 287 125 289 136
rect 294 125 296 136
rect 307 125 309 134
rect 329 129 331 135
rect 339 129 341 137
rect 346 129 348 137
rect 356 129 358 137
rect 363 129 365 137
rect 373 128 375 137
rect 396 128 398 137
rect 406 129 408 137
rect 413 129 415 137
rect 423 129 425 137
rect 430 129 432 137
rect 440 129 442 135
rect 463 128 465 137
rect 473 129 475 137
rect 480 129 482 137
rect 490 129 492 137
rect 497 129 499 137
rect 507 129 509 135
rect 529 123 531 132
rect 539 123 541 129
rect 549 123 551 129
rect 572 128 574 140
rect 579 128 581 140
rect 589 128 591 137
rect 599 128 601 137
rect 615 123 617 132
rect 13 22 15 31
rect 23 25 25 31
rect 33 25 35 31
rect 62 20 64 29
rect 75 18 77 29
rect 82 18 84 29
rect 102 22 104 31
rect 118 17 120 26
rect 128 17 130 26
rect 138 14 140 26
rect 145 14 147 26
rect 176 20 178 29
rect 189 18 191 29
rect 196 18 198 29
rect 216 22 218 31
rect 232 17 234 26
rect 242 17 244 26
rect 252 14 254 26
rect 259 14 261 26
rect 287 18 289 29
rect 294 18 296 29
rect 307 20 309 29
rect 329 19 331 25
rect 339 17 341 25
rect 346 17 348 25
rect 356 17 358 25
rect 363 17 365 25
rect 373 17 375 26
rect 396 17 398 26
rect 406 17 408 25
rect 413 17 415 25
rect 423 17 425 25
rect 430 17 432 25
rect 440 19 442 25
rect 463 17 465 26
rect 473 17 475 25
rect 480 17 482 25
rect 490 17 492 25
rect 497 17 499 25
rect 507 19 509 25
rect 529 22 531 31
rect 539 25 541 31
rect 549 25 551 31
rect 572 14 574 26
rect 579 14 581 26
rect 589 17 591 26
rect 599 17 601 26
rect 615 22 617 31
<< pmos >>
rect 13 237 15 255
rect 26 227 28 248
rect 33 227 35 248
rect 62 236 64 254
rect 72 234 74 247
rect 82 234 84 247
rect 110 227 112 254
rect 126 236 128 254
rect 136 236 138 254
rect 146 227 148 254
rect 176 236 178 254
rect 186 234 188 247
rect 196 234 198 247
rect 224 227 226 254
rect 240 236 242 254
rect 250 236 252 254
rect 260 227 262 254
rect 287 234 289 247
rect 297 234 299 247
rect 307 236 309 254
rect 329 247 331 255
rect 339 227 341 243
rect 346 227 348 243
rect 356 227 358 243
rect 363 227 365 243
rect 373 227 375 245
rect 396 227 398 245
rect 440 247 442 255
rect 406 227 408 243
rect 413 227 415 243
rect 423 227 425 243
rect 430 227 432 243
rect 463 227 465 245
rect 507 247 509 255
rect 473 227 475 243
rect 480 227 482 243
rect 490 227 492 243
rect 497 227 499 243
rect 529 237 531 255
rect 542 227 544 248
rect 549 227 551 248
rect 571 227 573 254
rect 581 236 583 254
rect 591 236 593 254
rect 607 227 609 254
rect 13 187 15 205
rect 26 194 28 215
rect 33 194 35 215
rect 62 188 64 206
rect 72 195 74 208
rect 82 195 84 208
rect 110 188 112 215
rect 126 188 128 206
rect 136 188 138 206
rect 146 188 148 215
rect 176 188 178 206
rect 186 195 188 208
rect 196 195 198 208
rect 224 188 226 215
rect 240 188 242 206
rect 250 188 252 206
rect 260 188 262 215
rect 287 195 289 208
rect 297 195 299 208
rect 307 188 309 206
rect 339 199 341 215
rect 346 199 348 215
rect 356 199 358 215
rect 363 199 365 215
rect 329 187 331 195
rect 373 197 375 215
rect 396 197 398 215
rect 406 199 408 215
rect 413 199 415 215
rect 423 199 425 215
rect 430 199 432 215
rect 463 197 465 215
rect 473 199 475 215
rect 480 199 482 215
rect 490 199 492 215
rect 497 199 499 215
rect 440 187 442 195
rect 507 187 509 195
rect 529 187 531 205
rect 542 194 544 215
rect 549 194 551 215
rect 571 188 573 215
rect 581 188 583 206
rect 591 188 593 206
rect 607 188 609 215
rect 13 93 15 111
rect 26 83 28 104
rect 33 83 35 104
rect 62 92 64 110
rect 72 90 74 103
rect 82 90 84 103
rect 110 83 112 110
rect 126 92 128 110
rect 136 92 138 110
rect 146 83 148 110
rect 176 92 178 110
rect 186 90 188 103
rect 196 90 198 103
rect 224 83 226 110
rect 240 92 242 110
rect 250 92 252 110
rect 260 83 262 110
rect 287 90 289 103
rect 297 90 299 103
rect 307 92 309 110
rect 329 103 331 111
rect 339 83 341 99
rect 346 83 348 99
rect 356 83 358 99
rect 363 83 365 99
rect 373 83 375 101
rect 396 83 398 101
rect 440 103 442 111
rect 406 83 408 99
rect 413 83 415 99
rect 423 83 425 99
rect 430 83 432 99
rect 463 83 465 101
rect 507 103 509 111
rect 473 83 475 99
rect 480 83 482 99
rect 490 83 492 99
rect 497 83 499 99
rect 529 93 531 111
rect 542 83 544 104
rect 549 83 551 104
rect 571 83 573 110
rect 581 92 583 110
rect 591 92 593 110
rect 607 83 609 110
rect 13 43 15 61
rect 26 50 28 71
rect 33 50 35 71
rect 62 44 64 62
rect 72 51 74 64
rect 82 51 84 64
rect 110 44 112 71
rect 126 44 128 62
rect 136 44 138 62
rect 146 44 148 71
rect 176 44 178 62
rect 186 51 188 64
rect 196 51 198 64
rect 224 44 226 71
rect 240 44 242 62
rect 250 44 252 62
rect 260 44 262 71
rect 287 51 289 64
rect 297 51 299 64
rect 307 44 309 62
rect 339 55 341 71
rect 346 55 348 71
rect 356 55 358 71
rect 363 55 365 71
rect 329 43 331 51
rect 373 53 375 71
rect 396 53 398 71
rect 406 55 408 71
rect 413 55 415 71
rect 423 55 425 71
rect 430 55 432 71
rect 463 53 465 71
rect 473 55 475 71
rect 480 55 482 71
rect 490 55 492 71
rect 497 55 499 71
rect 440 43 442 51
rect 507 43 509 51
rect 529 43 531 61
rect 542 50 544 71
rect 549 50 551 71
rect 571 44 573 71
rect 581 44 583 62
rect 591 44 593 62
rect 607 44 609 71
<< polyct0 >>
rect 15 260 17 262
rect 64 260 66 262
rect 134 260 136 262
rect 144 259 146 261
rect 178 260 180 262
rect 248 260 250 262
rect 258 259 260 261
rect 305 260 307 262
rect 354 266 356 268
rect 372 265 374 267
rect 397 265 399 267
rect 347 250 349 252
rect 415 266 417 268
rect 422 250 424 252
rect 464 265 466 267
rect 482 266 484 268
rect 489 250 491 252
rect 531 260 533 262
rect 573 259 575 261
rect 583 260 585 262
rect 15 180 17 182
rect 64 180 66 182
rect 134 180 136 182
rect 144 181 146 183
rect 178 180 180 182
rect 248 180 250 182
rect 258 181 260 183
rect 305 180 307 182
rect 347 190 349 192
rect 354 174 356 176
rect 422 190 424 192
rect 372 175 374 177
rect 397 175 399 177
rect 415 174 417 176
rect 489 190 491 192
rect 464 175 466 177
rect 482 174 484 176
rect 531 180 533 182
rect 573 181 575 183
rect 583 180 585 182
rect 15 116 17 118
rect 64 116 66 118
rect 134 116 136 118
rect 144 115 146 117
rect 178 116 180 118
rect 248 116 250 118
rect 258 115 260 117
rect 305 116 307 118
rect 354 122 356 124
rect 372 121 374 123
rect 397 121 399 123
rect 347 106 349 108
rect 415 122 417 124
rect 422 106 424 108
rect 464 121 466 123
rect 482 122 484 124
rect 489 106 491 108
rect 531 116 533 118
rect 573 115 575 117
rect 583 116 585 118
rect 15 36 17 38
rect 64 36 66 38
rect 134 36 136 38
rect 144 37 146 39
rect 178 36 180 38
rect 248 36 250 38
rect 258 37 260 39
rect 305 36 307 38
rect 347 46 349 48
rect 354 30 356 32
rect 422 46 424 48
rect 372 31 374 33
rect 397 31 399 33
rect 415 30 417 32
rect 489 46 491 48
rect 464 31 466 33
rect 482 30 484 32
rect 531 36 533 38
rect 573 37 575 39
rect 583 36 585 38
<< polyct1 >>
rect 25 260 27 262
rect 74 260 76 262
rect 35 253 37 255
rect 113 265 115 267
rect 84 252 86 254
rect 188 260 190 262
rect 97 252 99 254
rect 227 265 229 267
rect 198 252 200 254
rect 295 260 297 262
rect 211 252 213 254
rect 285 252 287 254
rect 337 260 339 262
rect 364 255 366 257
rect 405 255 407 257
rect 432 260 434 262
rect 324 240 326 242
rect 472 255 474 257
rect 499 260 501 262
rect 445 240 447 242
rect 541 260 543 262
rect 512 240 514 242
rect 604 265 606 267
rect 551 253 553 255
rect 620 252 622 254
rect 35 187 37 189
rect 25 180 27 182
rect 84 188 86 190
rect 97 188 99 190
rect 74 180 76 182
rect 198 188 200 190
rect 211 188 213 190
rect 285 188 287 190
rect 113 175 115 177
rect 188 180 190 182
rect 227 175 229 177
rect 324 200 326 202
rect 295 180 297 182
rect 445 200 447 202
rect 337 180 339 182
rect 364 185 366 187
rect 405 185 407 187
rect 512 200 514 202
rect 432 180 434 182
rect 472 185 474 187
rect 499 180 501 182
rect 551 187 553 189
rect 620 188 622 190
rect 541 180 543 182
rect 604 175 606 177
rect 25 116 27 118
rect 74 116 76 118
rect 35 109 37 111
rect 113 121 115 123
rect 84 108 86 110
rect 188 116 190 118
rect 97 108 99 110
rect 227 121 229 123
rect 198 108 200 110
rect 295 116 297 118
rect 211 108 213 110
rect 285 108 287 110
rect 337 116 339 118
rect 364 111 366 113
rect 405 111 407 113
rect 432 116 434 118
rect 324 96 326 98
rect 472 111 474 113
rect 499 116 501 118
rect 445 96 447 98
rect 541 116 543 118
rect 512 96 514 98
rect 604 121 606 123
rect 551 109 553 111
rect 620 108 622 110
rect 35 43 37 45
rect 25 36 27 38
rect 84 44 86 46
rect 97 44 99 46
rect 74 36 76 38
rect 198 44 200 46
rect 211 44 213 46
rect 285 44 287 46
rect 113 31 115 33
rect 188 36 190 38
rect 227 31 229 33
rect 324 56 326 58
rect 295 36 297 38
rect 445 56 447 58
rect 337 36 339 38
rect 364 41 366 43
rect 405 41 407 43
rect 512 56 514 58
rect 432 36 434 38
rect 472 41 474 43
rect 499 36 501 38
rect 551 43 553 45
rect 620 44 622 46
rect 541 36 543 38
rect 604 31 606 33
<< ndifct0 >>
rect 19 282 21 284
rect 38 282 40 284
rect 28 269 30 271
rect 87 276 89 278
rect 111 277 113 279
rect 97 269 99 271
rect 123 274 125 276
rect 201 276 203 278
rect 225 277 227 279
rect 211 269 213 271
rect 237 274 239 276
rect 282 276 284 278
rect 324 275 326 277
rect 334 275 336 277
rect 351 277 353 279
rect 368 277 370 279
rect 401 277 403 279
rect 418 277 420 279
rect 435 275 437 277
rect 445 275 447 277
rect 468 277 470 279
rect 485 277 487 279
rect 535 282 537 284
rect 502 275 504 277
rect 512 275 514 277
rect 554 282 556 284
rect 544 269 546 271
rect 594 274 596 276
rect 606 277 608 279
rect 620 269 622 271
rect 28 171 30 173
rect 19 158 21 160
rect 97 171 99 173
rect 87 164 89 166
rect 111 163 113 165
rect 38 158 40 160
rect 123 166 125 168
rect 211 171 213 173
rect 201 164 203 166
rect 225 163 227 165
rect 237 166 239 168
rect 282 164 284 166
rect 324 165 326 167
rect 334 165 336 167
rect 351 163 353 165
rect 368 163 370 165
rect 401 163 403 165
rect 418 163 420 165
rect 435 165 437 167
rect 445 165 447 167
rect 468 163 470 165
rect 485 163 487 165
rect 502 165 504 167
rect 512 165 514 167
rect 544 171 546 173
rect 535 158 537 160
rect 554 158 556 160
rect 594 166 596 168
rect 620 171 622 173
rect 606 163 608 165
rect 19 138 21 140
rect 38 138 40 140
rect 28 125 30 127
rect 87 132 89 134
rect 111 133 113 135
rect 97 125 99 127
rect 123 130 125 132
rect 201 132 203 134
rect 225 133 227 135
rect 211 125 213 127
rect 237 130 239 132
rect 282 132 284 134
rect 324 131 326 133
rect 334 131 336 133
rect 351 133 353 135
rect 368 133 370 135
rect 401 133 403 135
rect 418 133 420 135
rect 435 131 437 133
rect 445 131 447 133
rect 468 133 470 135
rect 485 133 487 135
rect 535 138 537 140
rect 502 131 504 133
rect 512 131 514 133
rect 554 138 556 140
rect 544 125 546 127
rect 594 130 596 132
rect 606 133 608 135
rect 620 125 622 127
rect 28 27 30 29
rect 19 14 21 16
rect 97 27 99 29
rect 87 20 89 22
rect 111 19 113 21
rect 38 14 40 16
rect 123 22 125 24
rect 211 27 213 29
rect 201 20 203 22
rect 225 19 227 21
rect 237 22 239 24
rect 282 20 284 22
rect 324 21 326 23
rect 334 21 336 23
rect 351 19 353 21
rect 368 19 370 21
rect 401 19 403 21
rect 418 19 420 21
rect 435 21 437 23
rect 445 21 447 23
rect 468 19 470 21
rect 485 19 487 21
rect 502 21 504 23
rect 512 21 514 23
rect 544 27 546 29
rect 535 14 537 16
rect 554 14 556 16
rect 594 22 596 24
rect 620 27 622 29
rect 606 19 608 21
<< ndifct1 >>
rect 68 286 70 288
rect 8 269 10 271
rect 151 286 153 288
rect 182 286 184 288
rect 57 274 59 276
rect 133 276 135 278
rect 265 286 267 288
rect 301 286 303 288
rect 171 274 173 276
rect 247 276 249 278
rect 312 274 314 276
rect 378 274 380 276
rect 391 274 393 276
rect 458 274 460 276
rect 566 286 568 288
rect 524 269 526 271
rect 584 276 586 278
rect 8 171 10 173
rect 57 166 59 168
rect 133 164 135 166
rect 68 154 70 156
rect 171 166 173 168
rect 151 154 153 156
rect 247 164 249 166
rect 182 154 184 156
rect 312 166 314 168
rect 265 154 267 156
rect 301 154 303 156
rect 378 166 380 168
rect 391 166 393 168
rect 458 166 460 168
rect 524 171 526 173
rect 584 164 586 166
rect 566 154 568 156
rect 68 142 70 144
rect 8 125 10 127
rect 151 142 153 144
rect 182 142 184 144
rect 57 130 59 132
rect 133 132 135 134
rect 265 142 267 144
rect 301 142 303 144
rect 171 130 173 132
rect 247 132 249 134
rect 312 130 314 132
rect 378 130 380 132
rect 391 130 393 132
rect 458 130 460 132
rect 566 142 568 144
rect 524 125 526 127
rect 584 132 586 134
rect 8 27 10 29
rect 57 22 59 24
rect 133 20 135 22
rect 68 10 70 12
rect 171 22 173 24
rect 151 10 153 12
rect 247 20 249 22
rect 182 10 184 12
rect 312 22 314 24
rect 265 10 267 12
rect 301 10 303 12
rect 378 22 380 24
rect 391 22 393 24
rect 458 22 460 24
rect 524 27 526 29
rect 584 20 586 22
rect 566 10 568 12
<< ntiect1 >>
rect 9 226 11 228
rect 58 226 60 228
rect 131 226 133 228
rect 172 226 174 228
rect 245 226 247 228
rect 311 226 313 228
rect 525 226 527 228
rect 586 226 588 228
rect 9 214 11 216
rect 58 214 60 216
rect 131 214 133 216
rect 172 214 174 216
rect 245 214 247 216
rect 311 214 313 216
rect 525 214 527 216
rect 586 214 588 216
rect 9 82 11 84
rect 58 82 60 84
rect 131 82 133 84
rect 172 82 174 84
rect 245 82 247 84
rect 311 82 313 84
rect 525 82 527 84
rect 586 82 588 84
rect 9 70 11 72
rect 58 70 60 72
rect 131 70 133 72
rect 172 70 174 72
rect 245 70 247 72
rect 311 70 313 72
rect 525 70 527 72
rect 586 70 588 72
<< ptiect1 >>
rect 9 286 11 288
rect 58 286 60 288
rect 98 286 100 288
rect 172 286 174 288
rect 212 286 214 288
rect 311 286 313 288
rect 525 286 527 288
rect 619 286 621 288
rect 9 154 11 156
rect 58 154 60 156
rect 98 154 100 156
rect 172 154 174 156
rect 212 154 214 156
rect 311 154 313 156
rect 525 154 527 156
rect 619 154 621 156
rect 9 142 11 144
rect 58 142 60 144
rect 98 142 100 144
rect 172 142 174 144
rect 212 142 214 144
rect 311 142 313 144
rect 525 142 527 144
rect 619 142 621 144
rect 9 10 11 12
rect 58 10 60 12
rect 98 10 100 12
rect 172 10 174 12
rect 212 10 214 12
rect 311 10 313 12
rect 525 10 527 12
rect 619 10 621 12
<< pdifct0 >>
rect 19 229 21 231
rect 38 236 40 238
rect 105 250 107 252
rect 67 238 69 240
rect 77 243 79 245
rect 77 236 79 238
rect 87 236 89 238
rect 115 236 117 238
rect 131 250 133 252
rect 131 243 133 245
rect 115 229 117 231
rect 151 235 153 237
rect 219 250 221 252
rect 181 238 183 240
rect 191 243 193 245
rect 191 236 193 238
rect 201 236 203 238
rect 229 236 231 238
rect 245 250 247 252
rect 245 243 247 245
rect 229 229 231 231
rect 265 235 267 237
rect 282 236 284 238
rect 292 243 294 245
rect 292 236 294 238
rect 302 238 304 240
rect 324 251 326 253
rect 334 229 336 231
rect 351 239 353 241
rect 368 229 370 231
rect 445 251 447 253
rect 401 229 403 231
rect 418 239 420 241
rect 435 229 437 231
rect 512 251 514 253
rect 468 229 470 231
rect 485 239 487 241
rect 502 229 504 231
rect 535 229 537 231
rect 554 236 556 238
rect 566 235 568 237
rect 586 250 588 252
rect 586 243 588 245
rect 602 236 604 238
rect 602 229 604 231
rect 612 250 614 252
rect 19 211 21 213
rect 38 204 40 206
rect 67 202 69 204
rect 77 204 79 206
rect 77 197 79 199
rect 87 204 89 206
rect 105 190 107 192
rect 115 211 117 213
rect 115 204 117 206
rect 131 197 133 199
rect 131 190 133 192
rect 151 205 153 207
rect 181 202 183 204
rect 191 204 193 206
rect 191 197 193 199
rect 201 204 203 206
rect 219 190 221 192
rect 229 211 231 213
rect 229 204 231 206
rect 245 197 247 199
rect 245 190 247 192
rect 334 211 336 213
rect 265 205 267 207
rect 282 204 284 206
rect 292 204 294 206
rect 292 197 294 199
rect 302 202 304 204
rect 351 201 353 203
rect 368 211 370 213
rect 324 189 326 191
rect 401 211 403 213
rect 418 201 420 203
rect 435 211 437 213
rect 468 211 470 213
rect 485 201 487 203
rect 502 211 504 213
rect 535 211 537 213
rect 445 189 447 191
rect 512 189 514 191
rect 554 204 556 206
rect 566 205 568 207
rect 602 211 604 213
rect 586 197 588 199
rect 586 190 588 192
rect 602 204 604 206
rect 612 190 614 192
rect 19 85 21 87
rect 38 92 40 94
rect 105 106 107 108
rect 67 94 69 96
rect 77 99 79 101
rect 77 92 79 94
rect 87 92 89 94
rect 115 92 117 94
rect 131 106 133 108
rect 131 99 133 101
rect 115 85 117 87
rect 151 91 153 93
rect 219 106 221 108
rect 181 94 183 96
rect 191 99 193 101
rect 191 92 193 94
rect 201 92 203 94
rect 229 92 231 94
rect 245 106 247 108
rect 245 99 247 101
rect 229 85 231 87
rect 265 91 267 93
rect 282 92 284 94
rect 292 99 294 101
rect 292 92 294 94
rect 302 94 304 96
rect 324 107 326 109
rect 334 85 336 87
rect 351 95 353 97
rect 368 85 370 87
rect 445 107 447 109
rect 401 85 403 87
rect 418 95 420 97
rect 435 85 437 87
rect 512 107 514 109
rect 468 85 470 87
rect 485 95 487 97
rect 502 85 504 87
rect 535 85 537 87
rect 554 92 556 94
rect 566 91 568 93
rect 586 106 588 108
rect 586 99 588 101
rect 602 92 604 94
rect 602 85 604 87
rect 612 106 614 108
rect 19 67 21 69
rect 38 60 40 62
rect 67 58 69 60
rect 77 60 79 62
rect 77 53 79 55
rect 87 60 89 62
rect 105 46 107 48
rect 115 67 117 69
rect 115 60 117 62
rect 131 53 133 55
rect 131 46 133 48
rect 151 61 153 63
rect 181 58 183 60
rect 191 60 193 62
rect 191 53 193 55
rect 201 60 203 62
rect 219 46 221 48
rect 229 67 231 69
rect 229 60 231 62
rect 245 53 247 55
rect 245 46 247 48
rect 334 67 336 69
rect 265 61 267 63
rect 282 60 284 62
rect 292 60 294 62
rect 292 53 294 55
rect 302 58 304 60
rect 351 57 353 59
rect 368 67 370 69
rect 324 45 326 47
rect 401 67 403 69
rect 418 57 420 59
rect 435 67 437 69
rect 468 67 470 69
rect 485 57 487 59
rect 502 67 504 69
rect 535 67 537 69
rect 445 45 447 47
rect 512 45 514 47
rect 554 60 556 62
rect 566 61 568 63
rect 602 67 604 69
rect 586 53 588 55
rect 586 46 588 48
rect 602 60 604 62
rect 612 46 614 48
<< pdifct1 >>
rect 8 246 10 248
rect 8 239 10 241
rect 57 250 59 252
rect 57 243 59 245
rect 141 243 143 245
rect 171 250 173 252
rect 171 243 173 245
rect 255 243 257 245
rect 312 250 314 252
rect 312 243 314 245
rect 378 236 380 238
rect 391 236 393 238
rect 458 236 460 238
rect 524 246 526 248
rect 524 239 526 241
rect 576 243 578 245
rect 8 201 10 203
rect 8 194 10 196
rect 57 197 59 199
rect 57 190 59 192
rect 141 197 143 199
rect 171 197 173 199
rect 171 190 173 192
rect 255 197 257 199
rect 312 197 314 199
rect 312 190 314 192
rect 378 204 380 206
rect 391 204 393 206
rect 458 204 460 206
rect 524 201 526 203
rect 524 194 526 196
rect 576 197 578 199
rect 8 102 10 104
rect 8 95 10 97
rect 57 106 59 108
rect 57 99 59 101
rect 141 99 143 101
rect 171 106 173 108
rect 171 99 173 101
rect 255 99 257 101
rect 312 106 314 108
rect 312 99 314 101
rect 378 92 380 94
rect 391 92 393 94
rect 458 92 460 94
rect 524 102 526 104
rect 524 95 526 97
rect 576 99 578 101
rect 8 57 10 59
rect 8 50 10 52
rect 57 53 59 55
rect 57 46 59 48
rect 141 53 143 55
rect 171 53 173 55
rect 171 46 173 48
rect 255 53 257 55
rect 312 53 314 55
rect 312 46 314 48
rect 378 60 380 62
rect 391 60 393 62
rect 458 60 460 62
rect 524 57 526 59
rect 524 50 526 52
rect 576 53 578 55
<< alu0 >>
rect 17 284 23 285
rect 17 282 19 284
rect 21 282 23 284
rect 17 281 23 282
rect 36 284 42 285
rect 36 282 38 284
rect 40 282 42 284
rect 36 281 42 282
rect 109 279 115 285
rect 71 278 91 279
rect 71 276 87 278
rect 89 276 91 278
rect 109 277 111 279
rect 113 277 115 279
rect 109 276 115 277
rect 122 276 126 278
rect 71 275 91 276
rect 14 271 32 272
rect 14 269 28 271
rect 30 269 32 271
rect 14 268 32 269
rect 14 262 18 268
rect 14 260 15 262
rect 17 260 18 262
rect 10 239 11 250
rect 14 247 18 260
rect 33 255 39 256
rect 59 272 60 274
rect 71 271 75 275
rect 122 274 123 276
rect 125 274 126 276
rect 63 267 75 271
rect 63 262 67 267
rect 63 260 64 262
rect 66 260 67 262
rect 14 243 29 247
rect 25 239 29 243
rect 63 248 67 260
rect 96 271 100 273
rect 96 269 97 271
rect 99 269 100 271
rect 96 263 100 269
rect 122 271 126 274
rect 122 267 146 271
rect 96 259 107 263
rect 63 245 80 248
rect 63 244 77 245
rect 76 243 77 244
rect 79 243 80 245
rect 65 240 71 241
rect 25 238 42 239
rect 25 236 38 238
rect 40 236 42 238
rect 25 235 42 236
rect 65 238 67 240
rect 69 238 71 240
rect 17 231 23 232
rect 17 229 19 231
rect 21 229 23 231
rect 65 229 71 238
rect 76 238 80 243
rect 103 253 107 259
rect 142 263 146 267
rect 122 262 138 263
rect 122 260 134 262
rect 136 260 138 262
rect 122 259 138 260
rect 142 261 147 263
rect 142 259 144 261
rect 146 259 147 261
rect 122 253 126 259
rect 142 257 147 259
rect 142 255 146 257
rect 103 252 126 253
rect 103 250 105 252
rect 107 250 126 252
rect 103 249 126 250
rect 76 236 77 238
rect 79 236 80 238
rect 76 234 80 236
rect 85 238 91 239
rect 85 236 87 238
rect 89 236 91 238
rect 85 229 91 236
rect 114 238 118 240
rect 114 236 115 238
rect 117 236 118 238
rect 114 231 118 236
rect 122 238 126 249
rect 130 252 146 255
rect 130 250 131 252
rect 133 251 146 252
rect 133 250 134 251
rect 130 245 134 250
rect 130 243 131 245
rect 133 243 134 245
rect 130 241 134 243
rect 223 279 229 285
rect 185 278 205 279
rect 185 276 201 278
rect 203 276 205 278
rect 223 277 225 279
rect 227 277 229 279
rect 223 276 229 277
rect 236 276 240 278
rect 185 275 205 276
rect 173 272 174 274
rect 185 271 189 275
rect 236 274 237 276
rect 239 274 240 276
rect 280 278 300 279
rect 280 276 282 278
rect 284 276 300 278
rect 280 275 300 276
rect 177 267 189 271
rect 177 262 181 267
rect 177 260 178 262
rect 180 260 181 262
rect 177 248 181 260
rect 210 271 214 273
rect 210 269 211 271
rect 213 269 214 271
rect 210 263 214 269
rect 236 271 240 274
rect 236 267 260 271
rect 210 259 221 263
rect 177 245 194 248
rect 177 244 191 245
rect 190 243 191 244
rect 193 243 194 245
rect 179 240 185 241
rect 179 238 181 240
rect 183 238 185 240
rect 122 237 155 238
rect 122 235 151 237
rect 153 235 155 237
rect 122 234 155 235
rect 114 229 115 231
rect 117 229 118 231
rect 179 229 185 238
rect 190 238 194 243
rect 217 253 221 259
rect 256 263 260 267
rect 236 262 252 263
rect 236 260 248 262
rect 250 260 252 262
rect 236 259 252 260
rect 256 261 261 263
rect 256 259 258 261
rect 260 259 261 261
rect 236 253 240 259
rect 256 257 261 259
rect 256 255 260 257
rect 217 252 240 253
rect 217 250 219 252
rect 221 250 240 252
rect 217 249 240 250
rect 190 236 191 238
rect 193 236 194 238
rect 190 234 194 236
rect 199 238 205 239
rect 199 236 201 238
rect 203 236 205 238
rect 199 229 205 236
rect 228 238 232 240
rect 228 236 229 238
rect 231 236 232 238
rect 228 231 232 236
rect 236 238 240 249
rect 244 252 260 255
rect 244 250 245 252
rect 247 251 260 252
rect 296 271 300 275
rect 311 272 312 274
rect 296 267 308 271
rect 304 262 308 267
rect 304 260 305 262
rect 307 260 308 262
rect 247 250 248 251
rect 244 245 248 250
rect 244 243 245 245
rect 247 243 248 245
rect 244 241 248 243
rect 304 248 308 260
rect 291 245 308 248
rect 291 243 292 245
rect 294 244 308 245
rect 322 277 328 278
rect 322 275 324 277
rect 326 275 328 277
rect 322 274 328 275
rect 332 277 338 285
rect 332 275 334 277
rect 336 275 338 277
rect 349 279 364 280
rect 349 277 351 279
rect 353 277 364 279
rect 349 276 364 277
rect 332 274 338 275
rect 322 254 326 274
rect 360 271 364 276
rect 367 279 371 285
rect 367 277 368 279
rect 370 277 371 279
rect 367 275 371 277
rect 346 268 357 270
rect 346 266 354 268
rect 356 266 357 268
rect 360 269 374 271
rect 360 267 375 269
rect 346 264 357 266
rect 370 265 372 267
rect 374 265 375 267
rect 346 254 350 264
rect 370 263 375 265
rect 322 253 350 254
rect 322 251 324 253
rect 326 252 350 253
rect 326 251 347 252
rect 322 250 347 251
rect 349 250 350 252
rect 366 253 367 259
rect 346 248 350 250
rect 294 243 295 244
rect 280 238 286 239
rect 236 237 269 238
rect 236 235 265 237
rect 267 235 269 237
rect 236 234 269 235
rect 280 236 282 238
rect 284 236 286 238
rect 228 229 229 231
rect 231 229 232 231
rect 280 229 286 236
rect 291 238 295 243
rect 370 246 374 263
rect 358 242 374 246
rect 291 236 292 238
rect 294 236 295 238
rect 291 234 295 236
rect 300 240 306 241
rect 300 238 302 240
rect 304 238 306 240
rect 300 229 306 238
rect 349 241 362 242
rect 349 239 351 241
rect 353 239 362 241
rect 349 238 362 239
rect 400 279 404 285
rect 400 277 401 279
rect 403 277 404 279
rect 400 275 404 277
rect 407 279 422 280
rect 407 277 418 279
rect 420 277 422 279
rect 407 276 422 277
rect 433 277 439 285
rect 467 279 471 285
rect 407 271 411 276
rect 433 275 435 277
rect 437 275 439 277
rect 433 274 439 275
rect 443 277 449 278
rect 443 275 445 277
rect 447 275 449 277
rect 443 274 449 275
rect 397 269 411 271
rect 396 267 411 269
rect 414 268 425 270
rect 396 265 397 267
rect 399 265 401 267
rect 396 263 401 265
rect 414 266 415 268
rect 417 266 425 268
rect 414 264 425 266
rect 397 246 401 263
rect 404 253 405 259
rect 421 254 425 264
rect 445 254 449 274
rect 421 253 449 254
rect 421 252 445 253
rect 421 250 422 252
rect 424 251 445 252
rect 447 251 449 253
rect 424 250 449 251
rect 467 277 468 279
rect 470 277 471 279
rect 467 275 471 277
rect 474 279 489 280
rect 474 277 485 279
rect 487 277 489 279
rect 474 276 489 277
rect 500 277 506 285
rect 533 284 539 285
rect 533 282 535 284
rect 537 282 539 284
rect 533 281 539 282
rect 552 284 558 285
rect 552 282 554 284
rect 556 282 558 284
rect 552 281 558 282
rect 604 279 610 285
rect 474 271 478 276
rect 500 275 502 277
rect 504 275 506 277
rect 500 274 506 275
rect 510 277 516 278
rect 510 275 512 277
rect 514 275 516 277
rect 510 274 516 275
rect 464 269 478 271
rect 421 248 425 250
rect 397 242 413 246
rect 409 241 422 242
rect 409 239 418 241
rect 420 239 422 241
rect 409 238 422 239
rect 463 267 478 269
rect 481 268 492 270
rect 463 265 464 267
rect 466 265 468 267
rect 463 263 468 265
rect 481 266 482 268
rect 484 266 492 268
rect 481 264 492 266
rect 464 246 468 263
rect 471 253 472 259
rect 488 254 492 264
rect 512 254 516 274
rect 593 276 597 278
rect 604 277 606 279
rect 608 277 610 279
rect 604 276 610 277
rect 488 253 516 254
rect 488 252 512 253
rect 488 250 489 252
rect 491 251 512 252
rect 514 251 516 253
rect 491 250 516 251
rect 530 271 548 272
rect 530 269 544 271
rect 546 269 548 271
rect 530 268 548 269
rect 488 248 492 250
rect 530 262 534 268
rect 530 260 531 262
rect 533 260 534 262
rect 464 242 480 246
rect 476 241 489 242
rect 476 239 485 241
rect 487 239 489 241
rect 476 238 489 239
rect 526 239 527 250
rect 530 247 534 260
rect 593 274 594 276
rect 596 274 597 276
rect 593 271 597 274
rect 549 255 555 256
rect 530 243 545 247
rect 541 239 545 243
rect 573 267 597 271
rect 573 263 577 267
rect 619 271 623 273
rect 619 269 620 271
rect 622 269 623 271
rect 572 261 577 263
rect 572 259 573 261
rect 575 259 577 261
rect 581 262 597 263
rect 581 260 583 262
rect 585 260 597 262
rect 581 259 597 260
rect 572 257 577 259
rect 573 255 577 257
rect 573 252 589 255
rect 573 251 586 252
rect 585 250 586 251
rect 588 250 589 252
rect 585 245 589 250
rect 585 243 586 245
rect 588 243 589 245
rect 585 241 589 243
rect 593 253 597 259
rect 619 263 623 269
rect 612 259 623 263
rect 612 253 616 259
rect 593 252 616 253
rect 593 250 612 252
rect 614 250 616 252
rect 593 249 616 250
rect 541 238 558 239
rect 593 238 597 249
rect 541 236 554 238
rect 556 236 558 238
rect 541 235 558 236
rect 564 237 597 238
rect 564 235 566 237
rect 568 235 597 237
rect 564 234 597 235
rect 601 238 605 240
rect 601 236 602 238
rect 604 236 605 238
rect 333 231 337 233
rect 333 229 334 231
rect 336 229 337 231
rect 366 231 372 232
rect 366 229 368 231
rect 370 229 372 231
rect 399 231 405 232
rect 399 229 401 231
rect 403 229 405 231
rect 434 231 438 233
rect 434 229 435 231
rect 437 229 438 231
rect 466 231 472 232
rect 466 229 468 231
rect 470 229 472 231
rect 501 231 505 233
rect 501 229 502 231
rect 504 229 505 231
rect 533 231 539 232
rect 533 229 535 231
rect 537 229 539 231
rect 601 231 605 236
rect 601 229 602 231
rect 604 229 605 231
rect 17 211 19 213
rect 21 211 23 213
rect 17 210 23 211
rect 25 206 42 207
rect 25 204 38 206
rect 40 204 42 206
rect 25 203 42 204
rect 65 204 71 213
rect 10 192 11 203
rect 25 199 29 203
rect 65 202 67 204
rect 69 202 71 204
rect 65 201 71 202
rect 76 206 80 208
rect 76 204 77 206
rect 79 204 80 206
rect 14 195 29 199
rect 76 199 80 204
rect 85 206 91 213
rect 114 211 115 213
rect 117 211 118 213
rect 85 204 87 206
rect 89 204 91 206
rect 85 203 91 204
rect 114 206 118 211
rect 114 204 115 206
rect 117 204 118 206
rect 114 202 118 204
rect 122 207 155 208
rect 122 205 151 207
rect 153 205 155 207
rect 122 204 155 205
rect 179 204 185 213
rect 76 198 77 199
rect 14 182 18 195
rect 63 197 77 198
rect 79 197 80 199
rect 63 194 80 197
rect 33 186 39 187
rect 14 180 15 182
rect 17 180 18 182
rect 14 174 18 180
rect 14 173 32 174
rect 14 171 28 173
rect 30 171 32 173
rect 14 170 32 171
rect 63 182 67 194
rect 122 193 126 204
rect 179 202 181 204
rect 183 202 185 204
rect 179 201 185 202
rect 190 206 194 208
rect 190 204 191 206
rect 193 204 194 206
rect 103 192 126 193
rect 103 190 105 192
rect 107 190 126 192
rect 103 189 126 190
rect 103 183 107 189
rect 63 180 64 182
rect 66 180 67 182
rect 63 175 67 180
rect 63 171 75 175
rect 59 168 60 170
rect 71 167 75 171
rect 96 179 107 183
rect 96 173 100 179
rect 122 183 126 189
rect 130 199 134 201
rect 130 197 131 199
rect 133 197 134 199
rect 130 192 134 197
rect 130 190 131 192
rect 133 191 134 192
rect 133 190 146 191
rect 130 187 146 190
rect 142 185 146 187
rect 142 183 147 185
rect 122 182 138 183
rect 122 180 134 182
rect 136 180 138 182
rect 122 179 138 180
rect 142 181 144 183
rect 146 181 147 183
rect 142 179 147 181
rect 96 171 97 173
rect 99 171 100 173
rect 96 169 100 171
rect 142 175 146 179
rect 122 171 146 175
rect 122 168 126 171
rect 71 166 91 167
rect 122 166 123 168
rect 125 166 126 168
rect 71 164 87 166
rect 89 164 91 166
rect 71 163 91 164
rect 109 165 115 166
rect 109 163 111 165
rect 113 163 115 165
rect 122 164 126 166
rect 190 199 194 204
rect 199 206 205 213
rect 228 211 229 213
rect 231 211 232 213
rect 199 204 201 206
rect 203 204 205 206
rect 199 203 205 204
rect 228 206 232 211
rect 228 204 229 206
rect 231 204 232 206
rect 228 202 232 204
rect 236 207 269 208
rect 236 205 265 207
rect 267 205 269 207
rect 236 204 269 205
rect 280 206 286 213
rect 280 204 282 206
rect 284 204 286 206
rect 190 198 191 199
rect 177 197 191 198
rect 193 197 194 199
rect 177 194 194 197
rect 177 182 181 194
rect 236 193 240 204
rect 280 203 286 204
rect 291 206 295 208
rect 291 204 292 206
rect 294 204 295 206
rect 217 192 240 193
rect 217 190 219 192
rect 221 190 240 192
rect 217 189 240 190
rect 217 183 221 189
rect 177 180 178 182
rect 180 180 181 182
rect 177 175 181 180
rect 177 171 189 175
rect 173 168 174 170
rect 17 160 23 161
rect 17 158 19 160
rect 21 158 23 160
rect 17 157 23 158
rect 36 160 42 161
rect 36 158 38 160
rect 40 158 42 160
rect 36 157 42 158
rect 109 157 115 163
rect 185 167 189 171
rect 210 179 221 183
rect 210 173 214 179
rect 236 183 240 189
rect 244 199 248 201
rect 244 197 245 199
rect 247 197 248 199
rect 244 192 248 197
rect 244 190 245 192
rect 247 191 248 192
rect 247 190 260 191
rect 244 187 260 190
rect 256 185 260 187
rect 291 199 295 204
rect 300 204 306 213
rect 333 211 334 213
rect 336 211 337 213
rect 333 209 337 211
rect 366 211 368 213
rect 370 211 372 213
rect 366 210 372 211
rect 399 211 401 213
rect 403 211 405 213
rect 399 210 405 211
rect 434 211 435 213
rect 437 211 438 213
rect 434 209 438 211
rect 466 211 468 213
rect 470 211 472 213
rect 466 210 472 211
rect 501 211 502 213
rect 504 211 505 213
rect 501 209 505 211
rect 533 211 535 213
rect 537 211 539 213
rect 533 210 539 211
rect 601 211 602 213
rect 604 211 605 213
rect 300 202 302 204
rect 304 202 306 204
rect 300 201 306 202
rect 291 197 292 199
rect 294 198 295 199
rect 294 197 308 198
rect 291 194 308 197
rect 256 183 261 185
rect 236 182 252 183
rect 236 180 248 182
rect 250 180 252 182
rect 236 179 252 180
rect 256 181 258 183
rect 260 181 261 183
rect 256 179 261 181
rect 210 171 211 173
rect 213 171 214 173
rect 210 169 214 171
rect 256 175 260 179
rect 236 171 260 175
rect 236 168 240 171
rect 185 166 205 167
rect 236 166 237 168
rect 239 166 240 168
rect 304 182 308 194
rect 349 203 362 204
rect 349 201 351 203
rect 353 201 362 203
rect 349 200 362 201
rect 358 196 374 200
rect 346 192 350 194
rect 304 180 305 182
rect 307 180 308 182
rect 304 175 308 180
rect 296 171 308 175
rect 296 167 300 171
rect 311 168 312 170
rect 185 164 201 166
rect 203 164 205 166
rect 185 163 205 164
rect 223 165 229 166
rect 223 163 225 165
rect 227 163 229 165
rect 236 164 240 166
rect 280 166 300 167
rect 280 164 282 166
rect 284 164 300 166
rect 280 163 300 164
rect 223 157 229 163
rect 322 191 347 192
rect 322 189 324 191
rect 326 190 347 191
rect 349 190 350 192
rect 326 189 350 190
rect 322 188 350 189
rect 322 168 326 188
rect 346 178 350 188
rect 366 183 367 189
rect 370 179 374 196
rect 346 176 357 178
rect 346 174 354 176
rect 356 174 357 176
rect 370 177 375 179
rect 370 175 372 177
rect 374 175 375 177
rect 346 172 357 174
rect 360 173 375 175
rect 360 171 374 173
rect 322 167 328 168
rect 322 165 324 167
rect 326 165 328 167
rect 322 164 328 165
rect 332 167 338 168
rect 332 165 334 167
rect 336 165 338 167
rect 360 166 364 171
rect 332 157 338 165
rect 349 165 364 166
rect 349 163 351 165
rect 353 163 364 165
rect 349 162 364 163
rect 367 165 371 167
rect 367 163 368 165
rect 370 163 371 165
rect 367 157 371 163
rect 409 203 422 204
rect 409 201 418 203
rect 420 201 422 203
rect 409 200 422 201
rect 397 196 413 200
rect 397 179 401 196
rect 476 203 489 204
rect 421 192 425 194
rect 404 183 405 189
rect 421 190 422 192
rect 424 191 449 192
rect 424 190 445 191
rect 421 189 445 190
rect 447 189 449 191
rect 421 188 449 189
rect 396 177 401 179
rect 421 178 425 188
rect 396 175 397 177
rect 399 175 401 177
rect 414 176 425 178
rect 396 173 411 175
rect 397 171 411 173
rect 414 174 415 176
rect 417 174 425 176
rect 414 172 425 174
rect 400 165 404 167
rect 400 163 401 165
rect 403 163 404 165
rect 400 157 404 163
rect 407 166 411 171
rect 445 168 449 188
rect 433 167 439 168
rect 407 165 422 166
rect 407 163 418 165
rect 420 163 422 165
rect 407 162 422 163
rect 433 165 435 167
rect 437 165 439 167
rect 433 157 439 165
rect 443 167 449 168
rect 443 165 445 167
rect 447 165 449 167
rect 443 164 449 165
rect 476 201 485 203
rect 487 201 489 203
rect 476 200 489 201
rect 464 196 480 200
rect 464 179 468 196
rect 564 207 597 208
rect 541 206 558 207
rect 541 204 554 206
rect 556 204 558 206
rect 564 205 566 207
rect 568 205 597 207
rect 564 204 597 205
rect 541 203 558 204
rect 488 192 492 194
rect 471 183 472 189
rect 488 190 489 192
rect 491 191 516 192
rect 491 190 512 191
rect 488 189 512 190
rect 514 189 516 191
rect 488 188 516 189
rect 463 177 468 179
rect 488 178 492 188
rect 463 175 464 177
rect 466 175 468 177
rect 481 176 492 178
rect 463 173 478 175
rect 464 171 478 173
rect 481 174 482 176
rect 484 174 492 176
rect 481 172 492 174
rect 467 165 471 167
rect 467 163 468 165
rect 470 163 471 165
rect 467 157 471 163
rect 474 166 478 171
rect 512 168 516 188
rect 526 192 527 203
rect 541 199 545 203
rect 530 195 545 199
rect 530 182 534 195
rect 585 199 589 201
rect 585 197 586 199
rect 588 197 589 199
rect 549 186 555 187
rect 530 180 531 182
rect 533 180 534 182
rect 530 174 534 180
rect 530 173 548 174
rect 530 171 544 173
rect 546 171 548 173
rect 530 170 548 171
rect 585 192 589 197
rect 585 191 586 192
rect 573 190 586 191
rect 588 190 589 192
rect 573 187 589 190
rect 593 193 597 204
rect 601 206 605 211
rect 601 204 602 206
rect 604 204 605 206
rect 601 202 605 204
rect 593 192 616 193
rect 593 190 612 192
rect 614 190 616 192
rect 593 189 616 190
rect 573 185 577 187
rect 572 183 577 185
rect 593 183 597 189
rect 572 181 573 183
rect 575 181 577 183
rect 572 179 577 181
rect 581 182 597 183
rect 581 180 583 182
rect 585 180 597 182
rect 581 179 597 180
rect 500 167 506 168
rect 474 165 489 166
rect 474 163 485 165
rect 487 163 489 165
rect 474 162 489 163
rect 500 165 502 167
rect 504 165 506 167
rect 500 157 506 165
rect 510 167 516 168
rect 510 165 512 167
rect 514 165 516 167
rect 510 164 516 165
rect 573 175 577 179
rect 612 183 616 189
rect 612 179 623 183
rect 573 171 597 175
rect 593 168 597 171
rect 619 173 623 179
rect 619 171 620 173
rect 622 171 623 173
rect 619 169 623 171
rect 593 166 594 168
rect 596 166 597 168
rect 593 164 597 166
rect 604 165 610 166
rect 604 163 606 165
rect 608 163 610 165
rect 533 160 539 161
rect 533 158 535 160
rect 537 158 539 160
rect 533 157 539 158
rect 552 160 558 161
rect 552 158 554 160
rect 556 158 558 160
rect 552 157 558 158
rect 604 157 610 163
rect 17 140 23 141
rect 17 138 19 140
rect 21 138 23 140
rect 17 137 23 138
rect 36 140 42 141
rect 36 138 38 140
rect 40 138 42 140
rect 36 137 42 138
rect 109 135 115 141
rect 71 134 91 135
rect 71 132 87 134
rect 89 132 91 134
rect 109 133 111 135
rect 113 133 115 135
rect 109 132 115 133
rect 122 132 126 134
rect 71 131 91 132
rect 14 127 32 128
rect 14 125 28 127
rect 30 125 32 127
rect 14 124 32 125
rect 14 118 18 124
rect 14 116 15 118
rect 17 116 18 118
rect 10 95 11 106
rect 14 103 18 116
rect 33 111 39 112
rect 59 128 60 130
rect 71 127 75 131
rect 122 130 123 132
rect 125 130 126 132
rect 63 123 75 127
rect 63 118 67 123
rect 63 116 64 118
rect 66 116 67 118
rect 14 99 29 103
rect 25 95 29 99
rect 63 104 67 116
rect 96 127 100 129
rect 96 125 97 127
rect 99 125 100 127
rect 96 119 100 125
rect 122 127 126 130
rect 122 123 146 127
rect 96 115 107 119
rect 63 101 80 104
rect 63 100 77 101
rect 76 99 77 100
rect 79 99 80 101
rect 65 96 71 97
rect 25 94 42 95
rect 25 92 38 94
rect 40 92 42 94
rect 25 91 42 92
rect 65 94 67 96
rect 69 94 71 96
rect 17 87 23 88
rect 17 85 19 87
rect 21 85 23 87
rect 65 85 71 94
rect 76 94 80 99
rect 103 109 107 115
rect 142 119 146 123
rect 122 118 138 119
rect 122 116 134 118
rect 136 116 138 118
rect 122 115 138 116
rect 142 117 147 119
rect 142 115 144 117
rect 146 115 147 117
rect 122 109 126 115
rect 142 113 147 115
rect 142 111 146 113
rect 103 108 126 109
rect 103 106 105 108
rect 107 106 126 108
rect 103 105 126 106
rect 76 92 77 94
rect 79 92 80 94
rect 76 90 80 92
rect 85 94 91 95
rect 85 92 87 94
rect 89 92 91 94
rect 85 85 91 92
rect 114 94 118 96
rect 114 92 115 94
rect 117 92 118 94
rect 114 87 118 92
rect 122 94 126 105
rect 130 108 146 111
rect 130 106 131 108
rect 133 107 146 108
rect 133 106 134 107
rect 130 101 134 106
rect 130 99 131 101
rect 133 99 134 101
rect 130 97 134 99
rect 223 135 229 141
rect 185 134 205 135
rect 185 132 201 134
rect 203 132 205 134
rect 223 133 225 135
rect 227 133 229 135
rect 223 132 229 133
rect 236 132 240 134
rect 185 131 205 132
rect 173 128 174 130
rect 185 127 189 131
rect 236 130 237 132
rect 239 130 240 132
rect 280 134 300 135
rect 280 132 282 134
rect 284 132 300 134
rect 280 131 300 132
rect 177 123 189 127
rect 177 118 181 123
rect 177 116 178 118
rect 180 116 181 118
rect 177 104 181 116
rect 210 127 214 129
rect 210 125 211 127
rect 213 125 214 127
rect 210 119 214 125
rect 236 127 240 130
rect 236 123 260 127
rect 210 115 221 119
rect 177 101 194 104
rect 177 100 191 101
rect 190 99 191 100
rect 193 99 194 101
rect 179 96 185 97
rect 179 94 181 96
rect 183 94 185 96
rect 122 93 155 94
rect 122 91 151 93
rect 153 91 155 93
rect 122 90 155 91
rect 114 85 115 87
rect 117 85 118 87
rect 179 85 185 94
rect 190 94 194 99
rect 217 109 221 115
rect 256 119 260 123
rect 236 118 252 119
rect 236 116 248 118
rect 250 116 252 118
rect 236 115 252 116
rect 256 117 261 119
rect 256 115 258 117
rect 260 115 261 117
rect 236 109 240 115
rect 256 113 261 115
rect 256 111 260 113
rect 217 108 240 109
rect 217 106 219 108
rect 221 106 240 108
rect 217 105 240 106
rect 190 92 191 94
rect 193 92 194 94
rect 190 90 194 92
rect 199 94 205 95
rect 199 92 201 94
rect 203 92 205 94
rect 199 85 205 92
rect 228 94 232 96
rect 228 92 229 94
rect 231 92 232 94
rect 228 87 232 92
rect 236 94 240 105
rect 244 108 260 111
rect 244 106 245 108
rect 247 107 260 108
rect 296 127 300 131
rect 311 128 312 130
rect 296 123 308 127
rect 304 118 308 123
rect 304 116 305 118
rect 307 116 308 118
rect 247 106 248 107
rect 244 101 248 106
rect 244 99 245 101
rect 247 99 248 101
rect 244 97 248 99
rect 304 104 308 116
rect 291 101 308 104
rect 291 99 292 101
rect 294 100 308 101
rect 322 133 328 134
rect 322 131 324 133
rect 326 131 328 133
rect 322 130 328 131
rect 332 133 338 141
rect 332 131 334 133
rect 336 131 338 133
rect 349 135 364 136
rect 349 133 351 135
rect 353 133 364 135
rect 349 132 364 133
rect 332 130 338 131
rect 322 110 326 130
rect 360 127 364 132
rect 367 135 371 141
rect 367 133 368 135
rect 370 133 371 135
rect 367 131 371 133
rect 346 124 357 126
rect 346 122 354 124
rect 356 122 357 124
rect 360 125 374 127
rect 360 123 375 125
rect 346 120 357 122
rect 370 121 372 123
rect 374 121 375 123
rect 346 110 350 120
rect 370 119 375 121
rect 322 109 350 110
rect 322 107 324 109
rect 326 108 350 109
rect 326 107 347 108
rect 322 106 347 107
rect 349 106 350 108
rect 366 109 367 115
rect 346 104 350 106
rect 294 99 295 100
rect 280 94 286 95
rect 236 93 269 94
rect 236 91 265 93
rect 267 91 269 93
rect 236 90 269 91
rect 280 92 282 94
rect 284 92 286 94
rect 228 85 229 87
rect 231 85 232 87
rect 280 85 286 92
rect 291 94 295 99
rect 370 102 374 119
rect 358 98 374 102
rect 291 92 292 94
rect 294 92 295 94
rect 291 90 295 92
rect 300 96 306 97
rect 300 94 302 96
rect 304 94 306 96
rect 300 85 306 94
rect 349 97 362 98
rect 349 95 351 97
rect 353 95 362 97
rect 349 94 362 95
rect 400 135 404 141
rect 400 133 401 135
rect 403 133 404 135
rect 400 131 404 133
rect 407 135 422 136
rect 407 133 418 135
rect 420 133 422 135
rect 407 132 422 133
rect 433 133 439 141
rect 467 135 471 141
rect 407 127 411 132
rect 433 131 435 133
rect 437 131 439 133
rect 433 130 439 131
rect 443 133 449 134
rect 443 131 445 133
rect 447 131 449 133
rect 443 130 449 131
rect 397 125 411 127
rect 396 123 411 125
rect 414 124 425 126
rect 396 121 397 123
rect 399 121 401 123
rect 396 119 401 121
rect 414 122 415 124
rect 417 122 425 124
rect 414 120 425 122
rect 397 102 401 119
rect 404 109 405 115
rect 421 110 425 120
rect 445 110 449 130
rect 421 109 449 110
rect 421 108 445 109
rect 421 106 422 108
rect 424 107 445 108
rect 447 107 449 109
rect 424 106 449 107
rect 467 133 468 135
rect 470 133 471 135
rect 467 131 471 133
rect 474 135 489 136
rect 474 133 485 135
rect 487 133 489 135
rect 474 132 489 133
rect 500 133 506 141
rect 533 140 539 141
rect 533 138 535 140
rect 537 138 539 140
rect 533 137 539 138
rect 552 140 558 141
rect 552 138 554 140
rect 556 138 558 140
rect 552 137 558 138
rect 604 135 610 141
rect 474 127 478 132
rect 500 131 502 133
rect 504 131 506 133
rect 500 130 506 131
rect 510 133 516 134
rect 510 131 512 133
rect 514 131 516 133
rect 510 130 516 131
rect 464 125 478 127
rect 421 104 425 106
rect 397 98 413 102
rect 409 97 422 98
rect 409 95 418 97
rect 420 95 422 97
rect 409 94 422 95
rect 463 123 478 125
rect 481 124 492 126
rect 463 121 464 123
rect 466 121 468 123
rect 463 119 468 121
rect 481 122 482 124
rect 484 122 492 124
rect 481 120 492 122
rect 464 102 468 119
rect 471 109 472 115
rect 488 110 492 120
rect 512 110 516 130
rect 593 132 597 134
rect 604 133 606 135
rect 608 133 610 135
rect 604 132 610 133
rect 488 109 516 110
rect 488 108 512 109
rect 488 106 489 108
rect 491 107 512 108
rect 514 107 516 109
rect 491 106 516 107
rect 530 127 548 128
rect 530 125 544 127
rect 546 125 548 127
rect 530 124 548 125
rect 488 104 492 106
rect 530 118 534 124
rect 530 116 531 118
rect 533 116 534 118
rect 464 98 480 102
rect 476 97 489 98
rect 476 95 485 97
rect 487 95 489 97
rect 476 94 489 95
rect 526 95 527 106
rect 530 103 534 116
rect 593 130 594 132
rect 596 130 597 132
rect 593 127 597 130
rect 549 111 555 112
rect 530 99 545 103
rect 541 95 545 99
rect 573 123 597 127
rect 573 119 577 123
rect 619 127 623 129
rect 619 125 620 127
rect 622 125 623 127
rect 572 117 577 119
rect 572 115 573 117
rect 575 115 577 117
rect 581 118 597 119
rect 581 116 583 118
rect 585 116 597 118
rect 581 115 597 116
rect 572 113 577 115
rect 573 111 577 113
rect 573 108 589 111
rect 573 107 586 108
rect 585 106 586 107
rect 588 106 589 108
rect 585 101 589 106
rect 585 99 586 101
rect 588 99 589 101
rect 585 97 589 99
rect 593 109 597 115
rect 619 119 623 125
rect 612 115 623 119
rect 612 109 616 115
rect 593 108 616 109
rect 593 106 612 108
rect 614 106 616 108
rect 593 105 616 106
rect 541 94 558 95
rect 593 94 597 105
rect 541 92 554 94
rect 556 92 558 94
rect 541 91 558 92
rect 564 93 597 94
rect 564 91 566 93
rect 568 91 597 93
rect 564 90 597 91
rect 601 94 605 96
rect 601 92 602 94
rect 604 92 605 94
rect 333 87 337 89
rect 333 85 334 87
rect 336 85 337 87
rect 366 87 372 88
rect 366 85 368 87
rect 370 85 372 87
rect 399 87 405 88
rect 399 85 401 87
rect 403 85 405 87
rect 434 87 438 89
rect 434 85 435 87
rect 437 85 438 87
rect 466 87 472 88
rect 466 85 468 87
rect 470 85 472 87
rect 501 87 505 89
rect 501 85 502 87
rect 504 85 505 87
rect 533 87 539 88
rect 533 85 535 87
rect 537 85 539 87
rect 601 87 605 92
rect 601 85 602 87
rect 604 85 605 87
rect 17 67 19 69
rect 21 67 23 69
rect 17 66 23 67
rect 25 62 42 63
rect 25 60 38 62
rect 40 60 42 62
rect 25 59 42 60
rect 65 60 71 69
rect 10 48 11 59
rect 25 55 29 59
rect 65 58 67 60
rect 69 58 71 60
rect 65 57 71 58
rect 76 62 80 64
rect 76 60 77 62
rect 79 60 80 62
rect 14 51 29 55
rect 76 55 80 60
rect 85 62 91 69
rect 114 67 115 69
rect 117 67 118 69
rect 85 60 87 62
rect 89 60 91 62
rect 85 59 91 60
rect 114 62 118 67
rect 114 60 115 62
rect 117 60 118 62
rect 114 58 118 60
rect 122 63 155 64
rect 122 61 151 63
rect 153 61 155 63
rect 122 60 155 61
rect 179 60 185 69
rect 76 54 77 55
rect 14 38 18 51
rect 63 53 77 54
rect 79 53 80 55
rect 63 50 80 53
rect 33 42 39 43
rect 14 36 15 38
rect 17 36 18 38
rect 14 30 18 36
rect 14 29 32 30
rect 14 27 28 29
rect 30 27 32 29
rect 14 26 32 27
rect 63 38 67 50
rect 122 49 126 60
rect 179 58 181 60
rect 183 58 185 60
rect 179 57 185 58
rect 190 62 194 64
rect 190 60 191 62
rect 193 60 194 62
rect 103 48 126 49
rect 103 46 105 48
rect 107 46 126 48
rect 103 45 126 46
rect 103 39 107 45
rect 63 36 64 38
rect 66 36 67 38
rect 63 31 67 36
rect 63 27 75 31
rect 59 24 60 26
rect 71 23 75 27
rect 96 35 107 39
rect 96 29 100 35
rect 122 39 126 45
rect 130 55 134 57
rect 130 53 131 55
rect 133 53 134 55
rect 130 48 134 53
rect 130 46 131 48
rect 133 47 134 48
rect 133 46 146 47
rect 130 43 146 46
rect 142 41 146 43
rect 142 39 147 41
rect 122 38 138 39
rect 122 36 134 38
rect 136 36 138 38
rect 122 35 138 36
rect 142 37 144 39
rect 146 37 147 39
rect 142 35 147 37
rect 96 27 97 29
rect 99 27 100 29
rect 96 25 100 27
rect 142 31 146 35
rect 122 27 146 31
rect 122 24 126 27
rect 71 22 91 23
rect 122 22 123 24
rect 125 22 126 24
rect 71 20 87 22
rect 89 20 91 22
rect 71 19 91 20
rect 109 21 115 22
rect 109 19 111 21
rect 113 19 115 21
rect 122 20 126 22
rect 190 55 194 60
rect 199 62 205 69
rect 228 67 229 69
rect 231 67 232 69
rect 199 60 201 62
rect 203 60 205 62
rect 199 59 205 60
rect 228 62 232 67
rect 228 60 229 62
rect 231 60 232 62
rect 228 58 232 60
rect 236 63 269 64
rect 236 61 265 63
rect 267 61 269 63
rect 236 60 269 61
rect 280 62 286 69
rect 280 60 282 62
rect 284 60 286 62
rect 190 54 191 55
rect 177 53 191 54
rect 193 53 194 55
rect 177 50 194 53
rect 177 38 181 50
rect 236 49 240 60
rect 280 59 286 60
rect 291 62 295 64
rect 291 60 292 62
rect 294 60 295 62
rect 217 48 240 49
rect 217 46 219 48
rect 221 46 240 48
rect 217 45 240 46
rect 217 39 221 45
rect 177 36 178 38
rect 180 36 181 38
rect 177 31 181 36
rect 177 27 189 31
rect 173 24 174 26
rect 17 16 23 17
rect 17 14 19 16
rect 21 14 23 16
rect 17 13 23 14
rect 36 16 42 17
rect 36 14 38 16
rect 40 14 42 16
rect 36 13 42 14
rect 109 13 115 19
rect 185 23 189 27
rect 210 35 221 39
rect 210 29 214 35
rect 236 39 240 45
rect 244 55 248 57
rect 244 53 245 55
rect 247 53 248 55
rect 244 48 248 53
rect 244 46 245 48
rect 247 47 248 48
rect 247 46 260 47
rect 244 43 260 46
rect 256 41 260 43
rect 291 55 295 60
rect 300 60 306 69
rect 333 67 334 69
rect 336 67 337 69
rect 333 65 337 67
rect 366 67 368 69
rect 370 67 372 69
rect 366 66 372 67
rect 399 67 401 69
rect 403 67 405 69
rect 399 66 405 67
rect 434 67 435 69
rect 437 67 438 69
rect 434 65 438 67
rect 466 67 468 69
rect 470 67 472 69
rect 466 66 472 67
rect 501 67 502 69
rect 504 67 505 69
rect 501 65 505 67
rect 533 67 535 69
rect 537 67 539 69
rect 533 66 539 67
rect 601 67 602 69
rect 604 67 605 69
rect 300 58 302 60
rect 304 58 306 60
rect 300 57 306 58
rect 291 53 292 55
rect 294 54 295 55
rect 294 53 308 54
rect 291 50 308 53
rect 256 39 261 41
rect 236 38 252 39
rect 236 36 248 38
rect 250 36 252 38
rect 236 35 252 36
rect 256 37 258 39
rect 260 37 261 39
rect 256 35 261 37
rect 210 27 211 29
rect 213 27 214 29
rect 210 25 214 27
rect 256 31 260 35
rect 236 27 260 31
rect 236 24 240 27
rect 185 22 205 23
rect 236 22 237 24
rect 239 22 240 24
rect 304 38 308 50
rect 349 59 362 60
rect 349 57 351 59
rect 353 57 362 59
rect 349 56 362 57
rect 358 52 374 56
rect 346 48 350 50
rect 304 36 305 38
rect 307 36 308 38
rect 304 31 308 36
rect 296 27 308 31
rect 296 23 300 27
rect 311 24 312 26
rect 185 20 201 22
rect 203 20 205 22
rect 185 19 205 20
rect 223 21 229 22
rect 223 19 225 21
rect 227 19 229 21
rect 236 20 240 22
rect 280 22 300 23
rect 280 20 282 22
rect 284 20 300 22
rect 280 19 300 20
rect 223 13 229 19
rect 322 47 347 48
rect 322 45 324 47
rect 326 46 347 47
rect 349 46 350 48
rect 326 45 350 46
rect 322 44 350 45
rect 322 24 326 44
rect 346 34 350 44
rect 366 39 367 45
rect 370 35 374 52
rect 346 32 357 34
rect 346 30 354 32
rect 356 30 357 32
rect 370 33 375 35
rect 370 31 372 33
rect 374 31 375 33
rect 346 28 357 30
rect 360 29 375 31
rect 360 27 374 29
rect 322 23 328 24
rect 322 21 324 23
rect 326 21 328 23
rect 322 20 328 21
rect 332 23 338 24
rect 332 21 334 23
rect 336 21 338 23
rect 360 22 364 27
rect 332 13 338 21
rect 349 21 364 22
rect 349 19 351 21
rect 353 19 364 21
rect 349 18 364 19
rect 367 21 371 23
rect 367 19 368 21
rect 370 19 371 21
rect 367 13 371 19
rect 409 59 422 60
rect 409 57 418 59
rect 420 57 422 59
rect 409 56 422 57
rect 397 52 413 56
rect 397 35 401 52
rect 476 59 489 60
rect 421 48 425 50
rect 404 39 405 45
rect 421 46 422 48
rect 424 47 449 48
rect 424 46 445 47
rect 421 45 445 46
rect 447 45 449 47
rect 421 44 449 45
rect 396 33 401 35
rect 421 34 425 44
rect 396 31 397 33
rect 399 31 401 33
rect 414 32 425 34
rect 396 29 411 31
rect 397 27 411 29
rect 414 30 415 32
rect 417 30 425 32
rect 414 28 425 30
rect 400 21 404 23
rect 400 19 401 21
rect 403 19 404 21
rect 400 13 404 19
rect 407 22 411 27
rect 445 24 449 44
rect 433 23 439 24
rect 407 21 422 22
rect 407 19 418 21
rect 420 19 422 21
rect 407 18 422 19
rect 433 21 435 23
rect 437 21 439 23
rect 433 13 439 21
rect 443 23 449 24
rect 443 21 445 23
rect 447 21 449 23
rect 443 20 449 21
rect 476 57 485 59
rect 487 57 489 59
rect 476 56 489 57
rect 464 52 480 56
rect 464 35 468 52
rect 564 63 597 64
rect 541 62 558 63
rect 541 60 554 62
rect 556 60 558 62
rect 564 61 566 63
rect 568 61 597 63
rect 564 60 597 61
rect 541 59 558 60
rect 488 48 492 50
rect 471 39 472 45
rect 488 46 489 48
rect 491 47 516 48
rect 491 46 512 47
rect 488 45 512 46
rect 514 45 516 47
rect 488 44 516 45
rect 463 33 468 35
rect 488 34 492 44
rect 463 31 464 33
rect 466 31 468 33
rect 481 32 492 34
rect 463 29 478 31
rect 464 27 478 29
rect 481 30 482 32
rect 484 30 492 32
rect 481 28 492 30
rect 467 21 471 23
rect 467 19 468 21
rect 470 19 471 21
rect 467 13 471 19
rect 474 22 478 27
rect 512 24 516 44
rect 526 48 527 59
rect 541 55 545 59
rect 530 51 545 55
rect 530 38 534 51
rect 585 55 589 57
rect 585 53 586 55
rect 588 53 589 55
rect 549 42 555 43
rect 530 36 531 38
rect 533 36 534 38
rect 530 30 534 36
rect 530 29 548 30
rect 530 27 544 29
rect 546 27 548 29
rect 530 26 548 27
rect 585 48 589 53
rect 585 47 586 48
rect 573 46 586 47
rect 588 46 589 48
rect 573 43 589 46
rect 593 49 597 60
rect 601 62 605 67
rect 601 60 602 62
rect 604 60 605 62
rect 601 58 605 60
rect 593 48 616 49
rect 593 46 612 48
rect 614 46 616 48
rect 593 45 616 46
rect 573 41 577 43
rect 572 39 577 41
rect 593 39 597 45
rect 572 37 573 39
rect 575 37 577 39
rect 572 35 577 37
rect 581 38 597 39
rect 581 36 583 38
rect 585 36 597 38
rect 581 35 597 36
rect 500 23 506 24
rect 474 21 489 22
rect 474 19 485 21
rect 487 19 489 21
rect 474 18 489 19
rect 500 21 502 23
rect 504 21 506 23
rect 500 13 506 21
rect 510 23 516 24
rect 510 21 512 23
rect 514 21 516 23
rect 510 20 516 21
rect 573 31 577 35
rect 612 39 616 45
rect 612 35 623 39
rect 573 27 597 31
rect 593 24 597 27
rect 619 29 623 35
rect 619 27 620 29
rect 622 27 623 29
rect 619 25 623 27
rect 593 22 594 24
rect 596 22 597 24
rect 593 20 597 22
rect 604 21 610 22
rect 604 19 606 21
rect 608 19 610 21
rect 533 16 539 17
rect 533 14 535 16
rect 537 14 539 16
rect 533 13 539 14
rect 552 16 558 17
rect 552 14 554 16
rect 556 14 558 16
rect 552 13 558 14
rect 604 13 610 19
<< via1 >>
rect 39 260 41 262
rect 80 269 82 271
rect 105 269 107 271
rect 88 245 90 247
rect 152 268 154 270
rect 97 245 99 247
rect 170 260 172 262
rect 194 269 196 271
rect 219 269 221 271
rect 202 245 204 247
rect 211 245 213 247
rect 266 253 268 255
rect 313 268 315 270
rect 330 268 332 270
rect 355 252 357 254
rect 332 244 334 246
rect 379 260 381 262
rect 406 260 408 262
rect 437 268 439 270
rect 457 268 459 270
rect 480 253 482 255
rect 505 268 507 270
rect 523 252 525 254
rect 504 244 506 246
rect 565 268 567 270
rect 88 195 90 197
rect 39 180 41 182
rect 97 195 99 197
rect 80 171 82 173
rect 105 171 107 173
rect 152 172 154 174
rect 202 195 204 197
rect 170 180 172 182
rect 211 195 213 197
rect 194 171 196 173
rect 266 187 268 189
rect 219 171 221 173
rect 332 196 334 198
rect 313 172 315 174
rect 330 172 332 174
rect 355 188 357 190
rect 379 180 381 182
rect 406 180 408 182
rect 437 172 439 174
rect 504 196 506 198
rect 480 187 482 189
rect 457 172 459 174
rect 505 172 507 174
rect 523 188 525 190
rect 565 172 567 174
rect 39 116 41 118
rect 80 125 82 127
rect 105 125 107 127
rect 88 101 90 103
rect 152 124 154 126
rect 97 101 99 103
rect 170 116 172 118
rect 194 125 196 127
rect 219 125 221 127
rect 202 101 204 103
rect 211 101 213 103
rect 266 109 268 111
rect 313 124 315 126
rect 330 124 332 126
rect 355 108 357 110
rect 332 100 334 102
rect 379 116 381 118
rect 406 116 408 118
rect 437 124 439 126
rect 457 124 459 126
rect 480 109 482 111
rect 505 124 507 126
rect 523 108 525 110
rect 504 100 506 102
rect 565 124 567 126
rect 88 51 90 53
rect 39 36 41 38
rect 97 51 99 53
rect 80 27 82 29
rect 105 27 107 29
rect 152 28 154 30
rect 202 51 204 53
rect 170 36 172 38
rect 211 51 213 53
rect 194 27 196 29
rect 266 43 268 45
rect 219 27 221 29
rect 332 52 334 54
rect 313 28 315 30
rect 330 28 332 30
rect 355 44 357 46
rect 379 36 381 38
rect 406 36 408 38
rect 437 28 439 30
rect 504 52 506 54
rect 480 43 482 45
rect 457 28 459 30
rect 505 28 507 30
rect 523 44 525 46
rect 565 28 567 30
<< labels >>
rlabel alu1 125 9 125 9 6 vss
rlabel alu1 125 73 125 73 6 vdd
rlabel alu1 73 73 73 73 6 vdd
rlabel alu1 73 9 73 9 6 vss
rlabel alu1 239 9 239 9 6 vss
rlabel alu1 239 73 239 73 6 vdd
rlabel alu1 187 73 187 73 6 vdd
rlabel alu1 187 9 187 9 6 vss
rlabel alu1 24 9 24 9 6 vss
rlabel alu1 24 73 24 73 6 vdd
rlabel via1 204 52 204 52 1 cin
rlabel alu1 298 9 298 9 4 vss
rlabel alu1 298 73 298 73 4 vdd
rlabel alu1 419 9 419 9 6 vss
rlabel alu1 419 73 419 73 6 vdd
rlabel alu1 352 9 352 9 4 vss
rlabel alu1 352 73 352 73 4 vdd
rlabel alu1 486 9 486 9 6 vss
rlabel alu1 486 73 486 73 6 vdd
rlabel via1 506 53 506 53 1 s1
rlabel alu1 514 61 514 61 1 s1
rlabel via1 332 53 332 53 1 s1
rlabel alu1 324 61 324 61 1 s1
rlabel alu1 447 61 447 61 1 s0
rlabel alu1 540 9 540 9 6 vss
rlabel alu1 540 73 540 73 6 vdd
rlabel alu1 594 9 594 9 4 vss
rlabel alu1 594 73 594 73 4 vdd
rlabel alu1 80 33 80 33 1 a0
rlabel via1 88 51 88 51 1 b0
rlabel alu1 282 53 282 53 1 b0
rlabel alu1 298 37 298 37 1 a0
rlabel alu1 540 37 540 37 1 a0
rlabel alu1 548 37 548 37 1 a0
rlabel alu1 540 45 540 45 1 b0
rlabel alu1 548 45 548 45 1 b0
rlabel alu1 556 53 556 53 1 b0
rlabel alu1 614 61 614 61 1 b0
rlabel alu1 622 53 622 53 1 b0
rlabel polyct1 606 33 606 33 1 a0
rlabel alu1 614 29 614 29 1 a0
rlabel alu1 290 33 290 33 1 a0
rlabel alu1 391 47 391 47 1 z0
rlabel alu1 399 61 399 61 1 z0
rlabel alu1 125 145 125 145 8 vss
rlabel alu1 125 81 125 81 8 vdd
rlabel alu1 73 81 73 81 8 vdd
rlabel alu1 73 145 73 145 8 vss
rlabel alu1 239 145 239 145 8 vss
rlabel alu1 239 81 239 81 8 vdd
rlabel alu1 187 81 187 81 8 vdd
rlabel alu1 187 145 187 145 8 vss
rlabel alu1 24 145 24 145 8 vss
rlabel alu1 24 81 24 81 8 vdd
rlabel alu1 298 145 298 145 2 vss
rlabel alu1 298 81 298 81 2 vdd
rlabel alu1 419 145 419 145 8 vss
rlabel alu1 419 81 419 81 8 vdd
rlabel alu1 352 145 352 145 2 vss
rlabel alu1 352 81 352 81 2 vdd
rlabel alu1 486 145 486 145 8 vss
rlabel alu1 486 81 486 81 8 vdd
rlabel via1 506 101 506 101 5 s1
rlabel alu1 514 93 514 93 5 s1
rlabel via1 332 101 332 101 5 s1
rlabel alu1 324 93 324 93 5 s1
rlabel alu1 447 93 447 93 5 s0
rlabel alu1 540 145 540 145 8 vss
rlabel alu1 540 81 540 81 8 vdd
rlabel alu1 594 145 594 145 2 vss
rlabel alu1 594 81 594 81 2 vdd
rlabel via1 204 102 204 102 1 cin1
rlabel alu1 8 39 8 39 1 cin1
rlabel alu1 80 121 80 121 1 a1
rlabel via1 88 103 88 103 1 b1
rlabel alu1 282 101 282 101 1 b1
rlabel alu1 290 121 290 121 1 a1
rlabel alu1 298 117 298 117 1 a1
rlabel alu1 391 107 391 107 1 z1
rlabel alu1 399 93 399 93 1 z1
rlabel alu1 540 117 540 117 1 a1
rlabel alu1 548 117 548 117 1 a1
rlabel alu1 540 109 540 109 1 b1
rlabel alu1 548 109 548 109 1 b1
rlabel alu1 556 101 556 101 1 b1
rlabel polyct1 606 121 606 121 1 a1
rlabel alu1 614 125 614 125 1 a1
rlabel alu1 622 101 622 101 1 b1
rlabel alu1 614 93 614 93 1 b1
rlabel alu1 8 115 8 115 1 cin2
rlabel alu1 125 153 125 153 6 vss
rlabel alu1 125 217 125 217 6 vdd
rlabel alu1 73 217 73 217 6 vdd
rlabel alu1 73 153 73 153 6 vss
rlabel alu1 239 153 239 153 6 vss
rlabel alu1 239 217 239 217 6 vdd
rlabel alu1 187 217 187 217 6 vdd
rlabel alu1 187 153 187 153 6 vss
rlabel alu1 24 153 24 153 6 vss
rlabel alu1 24 217 24 217 6 vdd
rlabel alu1 298 153 298 153 4 vss
rlabel alu1 298 217 298 217 4 vdd
rlabel alu1 419 153 419 153 6 vss
rlabel alu1 419 217 419 217 6 vdd
rlabel alu1 352 153 352 153 4 vss
rlabel alu1 352 217 352 217 4 vdd
rlabel alu1 486 153 486 153 6 vss
rlabel alu1 486 217 486 217 6 vdd
rlabel via1 506 197 506 197 1 s1
rlabel alu1 514 205 514 205 1 s1
rlabel via1 332 197 332 197 1 s1
rlabel alu1 324 205 324 205 1 s1
rlabel alu1 447 205 447 205 1 s0
rlabel alu1 540 153 540 153 6 vss
rlabel alu1 540 217 540 217 6 vdd
rlabel alu1 594 153 594 153 4 vss
rlabel alu1 594 217 594 217 4 vdd
rlabel alu1 125 289 125 289 8 vss
rlabel alu1 125 225 125 225 8 vdd
rlabel alu1 73 225 73 225 8 vdd
rlabel alu1 73 289 73 289 8 vss
rlabel alu1 239 289 239 289 8 vss
rlabel alu1 239 225 239 225 8 vdd
rlabel alu1 187 225 187 225 8 vdd
rlabel alu1 187 289 187 289 8 vss
rlabel alu1 24 289 24 289 8 vss
rlabel alu1 24 225 24 225 8 vdd
rlabel alu1 8 259 8 259 5 cout
rlabel alu1 298 289 298 289 2 vss
rlabel alu1 298 225 298 225 2 vdd
rlabel alu1 419 289 419 289 8 vss
rlabel alu1 419 225 419 225 8 vdd
rlabel alu1 352 289 352 289 2 vss
rlabel alu1 352 225 352 225 2 vdd
rlabel alu1 486 289 486 289 8 vss
rlabel alu1 486 225 486 225 8 vdd
rlabel via1 506 245 506 245 5 s1
rlabel alu1 514 237 514 237 5 s1
rlabel via1 332 245 332 245 5 s1
rlabel alu1 324 237 324 237 5 s1
rlabel alu1 447 237 447 237 5 s0
rlabel alu1 540 289 540 289 8 vss
rlabel alu1 540 225 540 225 8 vdd
rlabel alu1 594 289 594 289 2 vss
rlabel alu1 594 225 594 225 2 vdd
rlabel alu1 8 183 8 183 1 cin3
rlabel alu1 80 177 80 177 1 a2
rlabel via1 88 195 88 195 1 b2
rlabel alu1 282 197 282 197 1 b2
rlabel alu1 290 177 290 177 1 a2
rlabel alu1 298 181 298 181 1 a2
rlabel alu1 391 191 391 191 1 z2
rlabel alu1 399 205 399 205 1 z2
rlabel alu1 540 181 540 181 1 a2
rlabel alu1 548 181 548 181 1 a2
rlabel alu1 540 189 540 189 1 b2
rlabel alu1 548 189 548 189 1 b2
rlabel alu1 556 197 556 197 1 b2
rlabel alu1 614 205 614 205 1 b2
rlabel alu1 622 197 622 197 1 b2
rlabel polyct1 606 177 606 177 1 a2
rlabel alu1 614 173 614 173 1 a2
rlabel via1 204 196 204 196 1 cin2
rlabel via1 88 247 88 247 1 b3
rlabel alu1 80 265 80 265 1 a3
rlabel via1 204 246 204 246 1 cin3
rlabel alu1 282 245 282 245 1 b3
rlabel alu1 290 265 290 265 1 a3
rlabel alu1 298 261 298 261 1 a3
rlabel alu1 391 251 391 251 1 z3
rlabel alu1 399 237 399 237 1 z3
rlabel alu1 540 261 540 261 1 a3
rlabel alu1 548 261 548 261 1 a3
rlabel alu1 540 253 540 253 1 b3
rlabel alu1 548 253 548 253 1 b3
rlabel alu1 556 245 556 245 1 b3
rlabel polyct1 606 265 606 265 1 a3
rlabel alu1 614 269 614 269 1 a3
rlabel alu1 614 237 614 237 1 b3
rlabel alu1 622 245 622 245 1 b3
<< end >>
