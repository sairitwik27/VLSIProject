magic
tech scmos
timestamp 1607713436
<< ab >>
rect 4 5 44 77
rect 46 69 51 77
rect 53 69 157 77
rect 53 37 93 69
rect 94 37 157 69
rect 53 5 157 37
rect 167 69 271 77
rect 272 69 274 77
rect 167 37 207 69
rect 208 37 271 69
rect 167 5 271 37
rect 272 5 276 13
rect 278 5 318 77
rect 319 69 383 77
rect 322 13 383 69
rect 319 5 383 13
rect 387 5 451 77
rect 455 5 518 77
rect 520 69 560 77
rect 561 69 626 77
rect 627 69 632 77
rect 521 13 560 69
rect 563 13 626 69
rect 520 5 560 13
rect 562 5 632 13
rect 88 0 94 5
rect 202 0 208 5
<< nwell >>
rect -1 37 632 82
<< pwell >>
rect -1 0 632 37
<< poly >>
rect 26 71 28 75
rect 33 71 35 75
rect 13 61 15 66
rect 110 71 112 75
rect 62 62 64 66
rect 72 64 74 69
rect 82 64 84 69
rect 13 40 15 43
rect 26 40 28 50
rect 33 47 35 50
rect 33 45 39 47
rect 33 43 35 45
rect 37 43 39 45
rect 33 41 39 43
rect 13 38 19 40
rect 13 36 15 38
rect 17 36 19 38
rect 13 34 19 36
rect 23 38 29 40
rect 23 36 25 38
rect 27 36 29 38
rect 23 34 29 36
rect 13 31 15 34
rect 23 31 25 34
rect 33 31 35 41
rect 62 40 64 44
rect 72 40 74 51
rect 82 48 84 51
rect 82 46 88 48
rect 82 44 84 46
rect 86 44 88 46
rect 82 42 88 44
rect 95 46 101 48
rect 95 44 97 46
rect 99 44 101 46
rect 146 71 148 75
rect 126 62 128 66
rect 136 62 138 66
rect 224 71 226 75
rect 176 62 178 66
rect 186 64 188 69
rect 196 64 198 69
rect 95 42 101 44
rect 62 38 68 40
rect 62 36 64 38
rect 66 36 68 38
rect 62 34 68 36
rect 72 38 78 40
rect 72 36 74 38
rect 76 36 78 38
rect 72 34 78 36
rect 62 29 64 34
rect 75 29 77 34
rect 82 29 84 42
rect 99 41 101 42
rect 110 41 112 44
rect 126 41 128 44
rect 99 39 112 41
rect 118 39 128 41
rect 136 40 138 44
rect 146 41 148 44
rect 102 31 104 39
rect 118 35 120 39
rect 111 33 120 35
rect 132 38 138 40
rect 132 36 134 38
rect 136 36 138 38
rect 132 34 138 36
rect 142 39 148 41
rect 142 37 144 39
rect 146 37 148 39
rect 142 35 148 37
rect 176 40 178 44
rect 186 40 188 51
rect 196 48 198 51
rect 196 46 202 48
rect 196 44 198 46
rect 200 44 202 46
rect 196 42 202 44
rect 209 46 215 48
rect 209 44 211 46
rect 213 44 215 46
rect 260 71 262 75
rect 240 62 242 66
rect 250 62 252 66
rect 339 71 341 75
rect 346 71 348 75
rect 356 71 358 75
rect 363 71 365 75
rect 373 71 375 75
rect 396 71 398 75
rect 406 71 408 75
rect 413 71 415 75
rect 423 71 425 75
rect 430 71 432 75
rect 463 71 465 75
rect 473 71 475 75
rect 480 71 482 75
rect 490 71 492 75
rect 497 71 499 75
rect 287 64 289 69
rect 297 64 299 69
rect 307 62 309 66
rect 287 48 289 51
rect 283 46 289 48
rect 283 44 285 46
rect 287 44 289 46
rect 209 42 215 44
rect 176 38 182 40
rect 176 36 178 38
rect 180 36 182 38
rect 111 31 113 33
rect 115 31 120 33
rect 13 17 15 22
rect 23 20 25 25
rect 33 20 35 25
rect 62 16 64 20
rect 111 29 120 31
rect 136 31 138 34
rect 118 26 120 29
rect 128 26 130 30
rect 136 29 140 31
rect 138 26 140 29
rect 145 26 147 35
rect 176 34 182 36
rect 186 38 192 40
rect 186 36 188 38
rect 190 36 192 38
rect 186 34 192 36
rect 176 29 178 34
rect 189 29 191 34
rect 196 29 198 42
rect 213 41 215 42
rect 224 41 226 44
rect 240 41 242 44
rect 213 39 226 41
rect 232 39 242 41
rect 250 40 252 44
rect 260 41 262 44
rect 283 42 289 44
rect 216 31 218 39
rect 232 35 234 39
rect 225 33 234 35
rect 246 38 252 40
rect 246 36 248 38
rect 250 36 252 38
rect 246 34 252 36
rect 256 39 262 41
rect 256 37 258 39
rect 260 37 262 39
rect 256 35 262 37
rect 225 31 227 33
rect 229 31 234 33
rect 102 19 104 22
rect 75 13 77 18
rect 82 13 84 18
rect 102 17 107 19
rect 105 9 107 17
rect 118 13 120 17
rect 128 9 130 17
rect 176 16 178 20
rect 225 29 234 31
rect 250 31 252 34
rect 232 26 234 29
rect 242 26 244 30
rect 250 29 254 31
rect 252 26 254 29
rect 259 26 261 35
rect 287 29 289 42
rect 297 40 299 51
rect 322 58 328 60
rect 322 56 324 58
rect 326 56 328 58
rect 322 54 331 56
rect 329 51 331 54
rect 307 40 309 44
rect 293 38 299 40
rect 293 36 295 38
rect 297 36 299 38
rect 293 34 299 36
rect 303 38 309 40
rect 303 36 305 38
rect 307 36 309 38
rect 303 34 309 36
rect 294 29 296 34
rect 307 29 309 34
rect 216 19 218 22
rect 138 9 140 14
rect 145 9 147 14
rect 105 7 130 9
rect 189 13 191 18
rect 196 13 198 18
rect 216 17 221 19
rect 219 9 221 17
rect 232 13 234 17
rect 242 9 244 17
rect 329 25 331 43
rect 339 40 341 55
rect 346 50 348 55
rect 345 48 351 50
rect 345 46 347 48
rect 349 46 351 48
rect 345 44 351 46
rect 356 40 358 55
rect 363 45 365 55
rect 443 58 449 60
rect 443 56 445 58
rect 447 56 449 58
rect 335 38 341 40
rect 335 36 337 38
rect 339 36 341 38
rect 335 34 341 36
rect 339 25 341 34
rect 346 38 358 40
rect 362 43 368 45
rect 362 41 364 43
rect 366 41 368 43
rect 362 39 368 41
rect 346 25 348 38
rect 352 32 358 34
rect 352 30 354 32
rect 356 30 358 32
rect 352 28 358 30
rect 356 25 358 28
rect 363 25 365 39
rect 373 35 375 53
rect 396 35 398 53
rect 406 45 408 55
rect 403 43 409 45
rect 403 41 405 43
rect 407 41 409 43
rect 403 39 409 41
rect 413 40 415 55
rect 423 50 425 55
rect 420 48 426 50
rect 420 46 422 48
rect 424 46 426 48
rect 420 44 426 46
rect 430 40 432 55
rect 440 54 449 56
rect 440 51 442 54
rect 542 71 544 75
rect 549 71 551 75
rect 571 71 573 75
rect 529 61 531 66
rect 510 58 516 60
rect 510 56 512 58
rect 514 56 516 58
rect 370 33 376 35
rect 370 31 372 33
rect 374 31 376 33
rect 370 29 376 31
rect 395 33 401 35
rect 395 31 397 33
rect 399 31 401 33
rect 395 29 401 31
rect 373 26 375 29
rect 396 26 398 29
rect 252 9 254 14
rect 259 9 261 14
rect 287 13 289 18
rect 294 13 296 18
rect 219 7 244 9
rect 307 16 309 20
rect 329 9 331 19
rect 406 25 408 39
rect 413 38 425 40
rect 413 32 419 34
rect 413 30 415 32
rect 417 30 419 32
rect 413 28 419 30
rect 413 25 415 28
rect 423 25 425 38
rect 430 38 436 40
rect 430 36 432 38
rect 434 36 436 38
rect 430 34 436 36
rect 430 25 432 34
rect 440 25 442 43
rect 463 35 465 53
rect 473 45 475 55
rect 470 43 476 45
rect 470 41 472 43
rect 474 41 476 43
rect 470 39 476 41
rect 480 40 482 55
rect 490 50 492 55
rect 487 48 493 50
rect 487 46 489 48
rect 491 46 493 48
rect 487 44 493 46
rect 497 40 499 55
rect 507 54 516 56
rect 507 51 509 54
rect 462 33 468 35
rect 462 31 464 33
rect 466 31 468 33
rect 462 29 468 31
rect 463 26 465 29
rect 339 13 341 17
rect 346 9 348 17
rect 356 12 358 17
rect 363 12 365 17
rect 373 12 375 17
rect 396 12 398 17
rect 406 12 408 17
rect 413 12 415 17
rect 329 7 348 9
rect 423 9 425 17
rect 430 13 432 17
rect 440 9 442 19
rect 473 25 475 39
rect 480 38 492 40
rect 480 32 486 34
rect 480 30 482 32
rect 484 30 486 32
rect 480 28 486 30
rect 480 25 482 28
rect 490 25 492 38
rect 497 38 503 40
rect 497 36 499 38
rect 501 36 503 38
rect 497 34 503 36
rect 497 25 499 34
rect 507 25 509 43
rect 529 40 531 43
rect 542 40 544 50
rect 549 47 551 50
rect 549 45 555 47
rect 549 43 551 45
rect 553 43 555 45
rect 607 71 609 75
rect 581 62 583 66
rect 591 62 593 66
rect 618 46 624 48
rect 618 44 620 46
rect 622 44 624 46
rect 549 41 555 43
rect 571 41 573 44
rect 529 38 535 40
rect 529 36 531 38
rect 533 36 535 38
rect 529 34 535 36
rect 539 38 545 40
rect 539 36 541 38
rect 543 36 545 38
rect 539 34 545 36
rect 529 31 531 34
rect 539 31 541 34
rect 549 31 551 41
rect 571 39 577 41
rect 571 37 573 39
rect 575 37 577 39
rect 571 35 577 37
rect 581 40 583 44
rect 591 41 593 44
rect 607 41 609 44
rect 618 42 624 44
rect 618 41 620 42
rect 581 38 587 40
rect 591 39 601 41
rect 607 39 620 41
rect 581 36 583 38
rect 585 36 587 38
rect 572 26 574 35
rect 581 34 587 36
rect 599 35 601 39
rect 581 31 583 34
rect 579 29 583 31
rect 599 33 608 35
rect 599 31 604 33
rect 606 31 608 33
rect 615 31 617 39
rect 579 26 581 29
rect 589 26 591 30
rect 599 29 608 31
rect 599 26 601 29
rect 463 12 465 17
rect 473 12 475 17
rect 480 12 482 17
rect 423 7 442 9
rect 490 9 492 17
rect 497 13 499 17
rect 507 9 509 19
rect 529 17 531 22
rect 539 20 541 25
rect 549 20 551 25
rect 490 7 509 9
rect 615 19 617 22
rect 612 17 617 19
rect 572 9 574 14
rect 579 9 581 14
rect 589 9 591 17
rect 599 13 601 17
rect 612 9 614 17
rect 589 7 614 9
<< ndif >>
rect 6 29 13 31
rect 6 27 8 29
rect 10 27 13 29
rect 6 25 13 27
rect 8 22 13 25
rect 15 25 23 31
rect 25 29 33 31
rect 25 27 28 29
rect 30 27 33 29
rect 25 25 33 27
rect 35 25 42 31
rect 95 29 102 31
rect 57 26 62 29
rect 15 22 21 25
rect 17 18 21 22
rect 37 18 42 25
rect 55 24 62 26
rect 55 22 57 24
rect 59 22 62 24
rect 55 20 62 22
rect 64 20 75 29
rect 17 16 23 18
rect 17 14 19 16
rect 21 14 23 16
rect 17 12 23 14
rect 36 16 42 18
rect 66 18 75 20
rect 77 18 82 29
rect 84 24 89 29
rect 95 27 97 29
rect 99 27 102 29
rect 95 25 102 27
rect 84 22 91 24
rect 97 22 102 25
rect 104 26 109 31
rect 209 29 216 31
rect 171 26 176 29
rect 104 22 118 26
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 109 21 118 22
rect 109 19 111 21
rect 113 19 118 21
rect 36 14 38 16
rect 40 14 42 16
rect 36 12 42 14
rect 66 12 73 18
rect 109 17 118 19
rect 120 24 128 26
rect 120 22 123 24
rect 125 22 128 24
rect 120 17 128 22
rect 130 22 138 26
rect 130 20 133 22
rect 135 20 138 22
rect 130 17 138 20
rect 66 10 68 12
rect 70 10 73 12
rect 66 8 73 10
rect 133 14 138 17
rect 140 14 145 26
rect 147 14 155 26
rect 169 24 176 26
rect 169 22 171 24
rect 173 22 176 24
rect 169 20 176 22
rect 178 20 189 29
rect 180 18 189 20
rect 191 18 196 29
rect 198 24 203 29
rect 209 27 211 29
rect 213 27 216 29
rect 209 25 216 27
rect 198 22 205 24
rect 211 22 216 25
rect 218 26 223 31
rect 218 22 232 26
rect 198 20 201 22
rect 203 20 205 22
rect 198 18 205 20
rect 223 21 232 22
rect 223 19 225 21
rect 227 19 232 21
rect 149 12 155 14
rect 149 10 151 12
rect 153 10 155 12
rect 149 8 155 10
rect 180 12 187 18
rect 223 17 232 19
rect 234 24 242 26
rect 234 22 237 24
rect 239 22 242 24
rect 234 17 242 22
rect 244 22 252 26
rect 244 20 247 22
rect 249 20 252 22
rect 244 17 252 20
rect 180 10 182 12
rect 184 10 187 12
rect 180 8 187 10
rect 247 14 252 17
rect 254 14 259 26
rect 261 14 269 26
rect 282 24 287 29
rect 280 22 287 24
rect 280 20 282 22
rect 284 20 287 22
rect 280 18 287 20
rect 289 18 294 29
rect 296 20 307 29
rect 309 26 314 29
rect 309 24 316 26
rect 368 25 373 26
rect 309 22 312 24
rect 314 22 316 24
rect 309 20 316 22
rect 322 23 329 25
rect 322 21 324 23
rect 326 21 329 23
rect 296 18 305 20
rect 263 12 269 14
rect 263 10 265 12
rect 267 10 269 12
rect 263 8 269 10
rect 298 12 305 18
rect 322 19 329 21
rect 331 23 339 25
rect 331 21 334 23
rect 336 21 339 23
rect 331 19 339 21
rect 298 10 301 12
rect 303 10 305 12
rect 298 8 305 10
rect 333 17 339 19
rect 341 17 346 25
rect 348 21 356 25
rect 348 19 351 21
rect 353 19 356 21
rect 348 17 356 19
rect 358 17 363 25
rect 365 21 373 25
rect 365 19 368 21
rect 370 19 373 21
rect 365 17 373 19
rect 375 24 382 26
rect 375 22 378 24
rect 380 22 382 24
rect 375 20 382 22
rect 389 24 396 26
rect 389 22 391 24
rect 393 22 396 24
rect 389 20 396 22
rect 375 17 380 20
rect 391 17 396 20
rect 398 25 403 26
rect 398 21 406 25
rect 398 19 401 21
rect 403 19 406 21
rect 398 17 406 19
rect 408 17 413 25
rect 415 21 423 25
rect 415 19 418 21
rect 420 19 423 21
rect 415 17 423 19
rect 425 17 430 25
rect 432 23 440 25
rect 432 21 435 23
rect 437 21 440 23
rect 432 19 440 21
rect 442 23 449 25
rect 442 21 445 23
rect 447 21 449 23
rect 442 19 449 21
rect 456 24 463 26
rect 456 22 458 24
rect 460 22 463 24
rect 456 20 463 22
rect 432 17 438 19
rect 458 17 463 20
rect 465 25 470 26
rect 522 29 529 31
rect 522 27 524 29
rect 526 27 529 29
rect 522 25 529 27
rect 465 21 473 25
rect 465 19 468 21
rect 470 19 473 21
rect 465 17 473 19
rect 475 17 480 25
rect 482 21 490 25
rect 482 19 485 21
rect 487 19 490 21
rect 482 17 490 19
rect 492 17 497 25
rect 499 23 507 25
rect 499 21 502 23
rect 504 21 507 23
rect 499 19 507 21
rect 509 23 516 25
rect 509 21 512 23
rect 514 21 516 23
rect 524 22 529 25
rect 531 25 539 31
rect 541 29 549 31
rect 541 27 544 29
rect 546 27 549 29
rect 541 25 549 27
rect 551 25 558 31
rect 610 26 615 31
rect 531 22 537 25
rect 509 19 516 21
rect 499 17 505 19
rect 533 18 537 22
rect 553 18 558 25
rect 533 16 539 18
rect 533 14 535 16
rect 537 14 539 16
rect 533 12 539 14
rect 552 16 558 18
rect 552 14 554 16
rect 556 14 558 16
rect 552 12 558 14
rect 564 14 572 26
rect 574 14 579 26
rect 581 22 589 26
rect 581 20 584 22
rect 586 20 589 22
rect 581 17 589 20
rect 591 24 599 26
rect 591 22 594 24
rect 596 22 599 24
rect 591 17 599 22
rect 601 22 615 26
rect 617 29 624 31
rect 617 27 620 29
rect 622 27 624 29
rect 617 25 624 27
rect 617 22 622 25
rect 601 21 610 22
rect 601 19 606 21
rect 608 19 610 21
rect 601 17 610 19
rect 581 14 586 17
rect 564 12 570 14
rect 564 10 566 12
rect 568 10 570 12
rect 564 8 570 10
<< pdif >>
rect 17 69 26 71
rect 17 67 19 69
rect 21 67 26 69
rect 17 61 26 67
rect 6 59 13 61
rect 6 57 8 59
rect 10 57 13 59
rect 6 52 13 57
rect 6 50 8 52
rect 10 50 13 52
rect 6 48 13 50
rect 8 43 13 48
rect 15 50 26 61
rect 28 50 33 71
rect 35 64 40 71
rect 35 62 42 64
rect 66 62 72 64
rect 35 60 38 62
rect 40 60 42 62
rect 35 58 42 60
rect 35 50 40 58
rect 57 57 62 62
rect 55 55 62 57
rect 55 53 57 55
rect 59 53 62 55
rect 15 43 23 50
rect 55 48 62 53
rect 55 46 57 48
rect 59 46 62 48
rect 55 44 62 46
rect 64 60 72 62
rect 64 58 67 60
rect 69 58 72 60
rect 64 51 72 58
rect 74 62 82 64
rect 74 60 77 62
rect 79 60 82 62
rect 74 55 82 60
rect 74 53 77 55
rect 79 53 82 55
rect 74 51 82 53
rect 84 62 91 64
rect 84 60 87 62
rect 89 60 91 62
rect 84 51 91 60
rect 64 44 70 51
rect 105 50 110 71
rect 103 48 110 50
rect 103 46 105 48
rect 107 46 110 48
rect 103 44 110 46
rect 112 69 124 71
rect 112 67 115 69
rect 117 67 124 69
rect 112 62 124 67
rect 141 62 146 71
rect 112 60 115 62
rect 117 60 126 62
rect 112 44 126 60
rect 128 55 136 62
rect 128 53 131 55
rect 133 53 136 55
rect 128 48 136 53
rect 128 46 131 48
rect 133 46 136 48
rect 128 44 136 46
rect 138 55 146 62
rect 138 53 141 55
rect 143 53 146 55
rect 138 44 146 53
rect 148 65 153 71
rect 148 63 155 65
rect 148 61 151 63
rect 153 61 155 63
rect 180 62 186 64
rect 148 59 155 61
rect 148 44 153 59
rect 171 57 176 62
rect 169 55 176 57
rect 169 53 171 55
rect 173 53 176 55
rect 169 48 176 53
rect 169 46 171 48
rect 173 46 176 48
rect 169 44 176 46
rect 178 60 186 62
rect 178 58 181 60
rect 183 58 186 60
rect 178 51 186 58
rect 188 62 196 64
rect 188 60 191 62
rect 193 60 196 62
rect 188 55 196 60
rect 188 53 191 55
rect 193 53 196 55
rect 188 51 196 53
rect 198 62 205 64
rect 198 60 201 62
rect 203 60 205 62
rect 198 51 205 60
rect 178 44 184 51
rect 219 50 224 71
rect 217 48 224 50
rect 217 46 219 48
rect 221 46 224 48
rect 217 44 224 46
rect 226 69 238 71
rect 226 67 229 69
rect 231 67 238 69
rect 226 62 238 67
rect 255 62 260 71
rect 226 60 229 62
rect 231 60 240 62
rect 226 44 240 60
rect 242 55 250 62
rect 242 53 245 55
rect 247 53 250 55
rect 242 48 250 53
rect 242 46 245 48
rect 247 46 250 48
rect 242 44 250 46
rect 252 55 260 62
rect 252 53 255 55
rect 257 53 260 55
rect 252 44 260 53
rect 262 65 267 71
rect 262 63 269 65
rect 332 69 339 71
rect 332 67 334 69
rect 336 67 339 69
rect 262 61 265 63
rect 267 61 269 63
rect 262 59 269 61
rect 280 62 287 64
rect 280 60 282 62
rect 284 60 287 62
rect 262 44 267 59
rect 280 51 287 60
rect 289 62 297 64
rect 289 60 292 62
rect 294 60 297 62
rect 289 55 297 60
rect 289 53 292 55
rect 294 53 297 55
rect 289 51 297 53
rect 299 62 305 64
rect 299 60 307 62
rect 299 58 302 60
rect 304 58 307 60
rect 299 51 307 58
rect 301 44 307 51
rect 309 57 314 62
rect 332 59 339 67
rect 309 55 316 57
rect 309 53 312 55
rect 314 53 316 55
rect 309 48 316 53
rect 333 55 339 59
rect 341 55 346 71
rect 348 59 356 71
rect 348 57 351 59
rect 353 57 356 59
rect 348 55 356 57
rect 358 55 363 71
rect 365 69 373 71
rect 365 67 368 69
rect 370 67 373 69
rect 365 55 373 67
rect 333 51 337 55
rect 324 49 329 51
rect 309 46 312 48
rect 314 46 316 48
rect 309 44 316 46
rect 322 47 329 49
rect 322 45 324 47
rect 326 45 329 47
rect 322 43 329 45
rect 331 43 337 51
rect 368 53 373 55
rect 375 64 380 71
rect 391 64 396 71
rect 375 62 382 64
rect 375 60 378 62
rect 380 60 382 62
rect 375 58 382 60
rect 389 62 396 64
rect 389 60 391 62
rect 393 60 396 62
rect 389 58 396 60
rect 375 53 380 58
rect 391 53 396 58
rect 398 69 406 71
rect 398 67 401 69
rect 403 67 406 69
rect 398 55 406 67
rect 408 55 413 71
rect 415 59 423 71
rect 415 57 418 59
rect 420 57 423 59
rect 415 55 423 57
rect 425 55 430 71
rect 432 69 439 71
rect 432 67 435 69
rect 437 67 439 69
rect 432 59 439 67
rect 458 64 463 71
rect 456 62 463 64
rect 456 60 458 62
rect 460 60 463 62
rect 432 55 438 59
rect 456 58 463 60
rect 398 53 403 55
rect 434 51 438 55
rect 458 53 463 58
rect 465 69 473 71
rect 465 67 468 69
rect 470 67 473 69
rect 465 55 473 67
rect 475 55 480 71
rect 482 59 490 71
rect 482 57 485 59
rect 487 57 490 59
rect 482 55 490 57
rect 492 55 497 71
rect 499 69 506 71
rect 499 67 502 69
rect 504 67 506 69
rect 533 69 542 71
rect 499 59 506 67
rect 533 67 535 69
rect 537 67 542 69
rect 533 61 542 67
rect 499 55 505 59
rect 465 53 470 55
rect 434 43 440 51
rect 442 49 447 51
rect 442 47 449 49
rect 442 45 445 47
rect 447 45 449 47
rect 442 43 449 45
rect 501 51 505 55
rect 522 59 529 61
rect 522 57 524 59
rect 526 57 529 59
rect 522 52 529 57
rect 501 43 507 51
rect 509 49 514 51
rect 522 50 524 52
rect 526 50 529 52
rect 509 47 516 49
rect 522 48 529 50
rect 509 45 512 47
rect 514 45 516 47
rect 509 43 516 45
rect 524 43 529 48
rect 531 50 542 61
rect 544 50 549 71
rect 551 64 556 71
rect 566 65 571 71
rect 551 62 558 64
rect 551 60 554 62
rect 556 60 558 62
rect 551 58 558 60
rect 564 63 571 65
rect 564 61 566 63
rect 568 61 571 63
rect 564 59 571 61
rect 551 50 556 58
rect 531 43 539 50
rect 566 44 571 59
rect 573 62 578 71
rect 595 69 607 71
rect 595 67 602 69
rect 604 67 607 69
rect 595 62 607 67
rect 573 55 581 62
rect 573 53 576 55
rect 578 53 581 55
rect 573 44 581 53
rect 583 55 591 62
rect 583 53 586 55
rect 588 53 591 55
rect 583 48 591 53
rect 583 46 586 48
rect 588 46 591 48
rect 583 44 591 46
rect 593 60 602 62
rect 604 60 607 62
rect 593 44 607 60
rect 609 50 614 71
rect 609 48 616 50
rect 609 46 612 48
rect 614 46 616 48
rect 609 44 616 46
<< alu1 >>
rect 2 72 632 77
rect 2 70 9 72
rect 11 70 58 72
rect 60 70 131 72
rect 133 70 172 72
rect 174 70 245 72
rect 247 70 311 72
rect 313 70 525 72
rect 527 70 586 72
rect 588 70 632 72
rect 2 69 632 70
rect 6 63 10 64
rect 6 59 19 63
rect 6 57 8 59
rect 6 52 10 57
rect 6 50 8 52
rect 6 31 10 50
rect 38 53 42 56
rect 55 55 60 57
rect 55 53 57 55
rect 59 53 60 55
rect 95 58 107 64
rect 38 49 60 53
rect 38 47 42 49
rect 21 45 42 47
rect 21 43 35 45
rect 37 43 42 45
rect 55 48 60 49
rect 55 46 57 48
rect 59 46 60 48
rect 55 44 60 46
rect 87 53 91 56
rect 87 51 88 53
rect 90 51 91 53
rect 6 29 11 31
rect 6 27 8 29
rect 10 27 11 29
rect 6 25 11 27
rect 21 38 42 39
rect 21 36 25 38
rect 27 36 39 38
rect 41 36 42 38
rect 21 35 42 36
rect 38 26 42 35
rect 55 24 59 44
rect 87 47 91 51
rect 78 46 91 47
rect 78 44 84 46
rect 86 44 91 46
rect 78 43 91 44
rect 95 53 100 58
rect 95 51 97 53
rect 99 51 100 53
rect 95 46 100 51
rect 95 44 97 46
rect 99 44 100 46
rect 95 42 100 44
rect 70 38 84 39
rect 70 36 74 38
rect 76 36 84 38
rect 70 35 84 36
rect 55 22 57 24
rect 59 22 67 24
rect 55 18 67 22
rect 79 29 84 35
rect 79 27 80 29
rect 82 27 84 29
rect 79 26 84 27
rect 111 33 116 40
rect 139 55 155 56
rect 139 53 141 55
rect 143 53 155 55
rect 139 51 155 53
rect 111 32 113 33
rect 103 31 113 32
rect 115 31 116 33
rect 103 29 116 31
rect 103 27 105 29
rect 107 27 116 29
rect 103 26 116 27
rect 151 30 155 51
rect 151 28 152 30
rect 154 28 155 30
rect 151 23 155 28
rect 131 22 155 23
rect 131 20 133 22
rect 135 20 155 22
rect 131 19 155 20
rect 169 55 174 57
rect 169 53 171 55
rect 173 53 174 55
rect 209 58 221 64
rect 169 48 174 53
rect 169 46 171 48
rect 173 46 174 48
rect 169 44 174 46
rect 201 53 205 56
rect 201 51 202 53
rect 204 51 205 53
rect 169 38 173 44
rect 169 36 170 38
rect 172 36 173 38
rect 169 24 173 36
rect 201 47 205 51
rect 192 46 205 47
rect 192 44 198 46
rect 200 44 205 46
rect 192 43 205 44
rect 209 53 214 58
rect 209 51 211 53
rect 213 51 214 53
rect 209 46 214 51
rect 209 44 211 46
rect 213 44 214 46
rect 209 42 214 44
rect 184 38 198 39
rect 184 36 188 38
rect 190 36 198 38
rect 184 35 198 36
rect 169 22 171 24
rect 173 22 181 24
rect 169 18 181 22
rect 193 29 198 35
rect 193 27 194 29
rect 196 27 198 29
rect 193 26 198 27
rect 225 33 230 40
rect 253 55 269 56
rect 253 53 255 55
rect 257 53 269 55
rect 253 51 269 53
rect 265 45 269 51
rect 265 43 266 45
rect 268 43 269 45
rect 280 47 284 56
rect 322 58 327 64
rect 369 62 382 63
rect 369 60 378 62
rect 380 60 382 62
rect 311 55 316 57
rect 280 46 293 47
rect 280 44 285 46
rect 287 44 293 46
rect 280 43 293 44
rect 225 32 227 33
rect 217 31 227 32
rect 229 31 230 33
rect 217 29 230 31
rect 217 27 219 29
rect 221 27 230 29
rect 217 26 230 27
rect 265 23 269 43
rect 287 38 301 39
rect 287 36 295 38
rect 297 36 301 38
rect 287 35 301 36
rect 311 53 312 55
rect 314 53 316 55
rect 311 48 316 53
rect 322 56 324 58
rect 326 56 327 58
rect 369 59 382 60
rect 322 55 327 56
rect 322 54 335 55
rect 322 52 332 54
rect 334 52 335 54
rect 322 51 335 52
rect 311 46 312 48
rect 314 46 316 48
rect 311 44 316 46
rect 287 26 292 35
rect 312 30 316 44
rect 312 28 313 30
rect 315 28 316 30
rect 312 24 316 28
rect 245 22 269 23
rect 245 20 247 22
rect 249 20 269 22
rect 245 19 269 20
rect 304 22 312 24
rect 314 22 316 24
rect 304 18 316 22
rect 336 38 342 40
rect 336 36 337 38
rect 339 36 342 38
rect 336 31 342 36
rect 329 30 342 31
rect 329 28 330 30
rect 332 28 342 30
rect 354 46 366 48
rect 354 44 355 46
rect 357 44 366 46
rect 354 43 366 44
rect 354 42 364 43
rect 362 41 364 42
rect 362 34 366 41
rect 378 38 382 59
rect 378 36 379 38
rect 381 36 382 38
rect 329 27 342 28
rect 378 26 382 36
rect 377 24 382 26
rect 377 22 378 24
rect 380 22 382 24
rect 377 20 382 22
rect 378 18 382 20
rect 389 62 402 63
rect 389 60 391 62
rect 393 60 402 62
rect 389 59 402 60
rect 389 26 393 59
rect 444 58 449 64
rect 444 56 445 58
rect 447 56 449 58
rect 444 55 449 56
rect 436 51 449 55
rect 456 62 469 63
rect 456 60 458 62
rect 460 60 469 62
rect 456 59 469 60
rect 405 43 417 48
rect 407 42 417 43
rect 407 41 409 42
rect 405 38 409 41
rect 405 36 406 38
rect 408 36 409 38
rect 405 34 409 36
rect 429 38 435 40
rect 429 36 432 38
rect 434 36 435 38
rect 429 31 435 36
rect 429 30 442 31
rect 429 28 437 30
rect 439 28 442 30
rect 429 27 442 28
rect 389 24 394 26
rect 389 22 391 24
rect 393 22 394 24
rect 389 20 394 22
rect 389 18 393 20
rect 456 30 460 59
rect 511 58 516 64
rect 511 56 512 58
rect 514 56 516 58
rect 511 55 516 56
rect 503 54 516 55
rect 503 52 504 54
rect 506 52 516 54
rect 503 51 516 52
rect 522 63 526 64
rect 522 59 535 63
rect 522 57 524 59
rect 522 52 526 57
rect 522 50 524 52
rect 472 45 484 48
rect 472 43 480 45
rect 482 43 484 45
rect 474 42 484 43
rect 474 41 476 42
rect 456 28 457 30
rect 459 28 460 30
rect 472 34 476 41
rect 456 26 460 28
rect 496 38 502 40
rect 496 36 499 38
rect 501 36 502 38
rect 496 31 502 36
rect 496 30 509 31
rect 496 28 505 30
rect 507 28 509 30
rect 496 27 509 28
rect 456 24 461 26
rect 456 22 458 24
rect 460 22 461 24
rect 456 20 461 22
rect 456 18 460 20
rect 522 46 526 50
rect 522 44 523 46
rect 525 44 526 46
rect 522 31 526 44
rect 554 47 558 56
rect 537 45 558 47
rect 537 43 551 45
rect 553 43 558 45
rect 564 55 580 56
rect 564 53 576 55
rect 578 53 580 55
rect 564 51 580 53
rect 522 29 527 31
rect 522 27 524 29
rect 526 27 527 29
rect 522 25 527 27
rect 537 38 558 39
rect 537 36 541 38
rect 543 36 558 38
rect 537 35 558 36
rect 554 26 558 35
rect 564 30 568 51
rect 612 58 624 64
rect 564 28 565 30
rect 567 28 568 30
rect 564 23 568 28
rect 603 33 608 40
rect 619 46 624 58
rect 619 44 620 46
rect 622 44 624 46
rect 619 42 624 44
rect 603 31 604 33
rect 606 32 608 33
rect 606 31 616 32
rect 603 26 616 31
rect 564 22 588 23
rect 564 20 584 22
rect 586 20 588 22
rect 564 19 588 20
rect 2 12 632 13
rect 2 10 9 12
rect 11 10 58 12
rect 60 10 68 12
rect 70 10 98 12
rect 100 10 151 12
rect 153 10 172 12
rect 174 10 182 12
rect 184 10 212 12
rect 214 10 265 12
rect 267 10 301 12
rect 303 10 311 12
rect 313 10 525 12
rect 527 10 566 12
rect 568 10 619 12
rect 621 10 632 12
rect 2 5 632 10
<< alu2 >>
rect 331 54 508 55
rect 87 53 100 54
rect 87 51 88 53
rect 90 51 97 53
rect 99 51 100 53
rect 87 50 100 51
rect 201 53 214 54
rect 201 51 202 53
rect 204 51 211 53
rect 213 51 214 53
rect 331 52 332 54
rect 334 52 504 54
rect 506 52 508 54
rect 331 51 508 52
rect 201 50 214 51
rect 265 46 359 47
rect 265 45 355 46
rect 265 43 266 45
rect 268 44 355 45
rect 357 44 359 46
rect 268 43 359 44
rect 265 42 359 43
rect 479 46 526 47
rect 479 45 523 46
rect 479 43 480 45
rect 482 44 523 45
rect 525 44 526 46
rect 482 43 526 44
rect 479 42 526 43
rect 38 38 173 39
rect 38 36 39 38
rect 41 36 170 38
rect 172 36 173 38
rect 38 35 173 36
rect 378 38 409 39
rect 378 36 379 38
rect 381 36 406 38
rect 408 36 409 38
rect 378 35 409 36
rect 79 29 111 31
rect 79 27 80 29
rect 82 27 105 29
rect 107 27 111 29
rect 79 26 111 27
rect 151 30 225 31
rect 151 28 152 30
rect 154 29 225 30
rect 154 28 194 29
rect 151 27 194 28
rect 196 27 219 29
rect 221 27 225 29
rect 312 30 333 31
rect 312 28 313 30
rect 315 28 330 30
rect 332 28 333 30
rect 312 27 333 28
rect 436 30 460 31
rect 436 28 437 30
rect 439 28 457 30
rect 459 28 460 30
rect 436 27 460 28
rect 504 30 568 31
rect 504 28 505 30
rect 507 28 565 30
rect 567 28 568 30
rect 504 27 568 28
rect 151 26 225 27
<< ptie >>
rect 7 12 13 14
rect 56 12 62 14
rect 7 10 9 12
rect 11 10 13 12
rect 7 8 13 10
rect 56 10 58 12
rect 60 10 62 12
rect 56 8 62 10
rect 96 12 102 14
rect 96 10 98 12
rect 100 10 102 12
rect 96 8 102 10
rect 170 12 176 14
rect 170 10 172 12
rect 174 10 176 12
rect 170 8 176 10
rect 210 12 216 14
rect 210 10 212 12
rect 214 10 216 12
rect 210 8 216 10
rect 309 12 315 14
rect 309 10 311 12
rect 313 10 315 12
rect 309 8 315 10
rect 523 12 529 14
rect 523 10 525 12
rect 527 10 529 12
rect 523 8 529 10
rect 617 12 623 14
rect 617 10 619 12
rect 621 10 623 12
rect 617 8 623 10
<< ntie >>
rect 7 72 13 74
rect 7 70 9 72
rect 11 70 13 72
rect 56 72 62 74
rect 7 68 13 70
rect 56 70 58 72
rect 60 70 62 72
rect 129 72 135 74
rect 56 68 62 70
rect 129 70 131 72
rect 133 70 135 72
rect 170 72 176 74
rect 129 68 135 70
rect 170 70 172 72
rect 174 70 176 72
rect 243 72 249 74
rect 170 68 176 70
rect 243 70 245 72
rect 247 70 249 72
rect 309 72 315 74
rect 243 68 249 70
rect 309 70 311 72
rect 313 70 315 72
rect 523 72 529 74
rect 309 68 315 70
rect 523 70 525 72
rect 527 70 529 72
rect 584 72 590 74
rect 523 68 529 70
rect 584 70 586 72
rect 588 70 590 72
rect 584 68 590 70
<< nmos >>
rect 13 22 15 31
rect 23 25 25 31
rect 33 25 35 31
rect 62 20 64 29
rect 75 18 77 29
rect 82 18 84 29
rect 102 22 104 31
rect 118 17 120 26
rect 128 17 130 26
rect 138 14 140 26
rect 145 14 147 26
rect 176 20 178 29
rect 189 18 191 29
rect 196 18 198 29
rect 216 22 218 31
rect 232 17 234 26
rect 242 17 244 26
rect 252 14 254 26
rect 259 14 261 26
rect 287 18 289 29
rect 294 18 296 29
rect 307 20 309 29
rect 329 19 331 25
rect 339 17 341 25
rect 346 17 348 25
rect 356 17 358 25
rect 363 17 365 25
rect 373 17 375 26
rect 396 17 398 26
rect 406 17 408 25
rect 413 17 415 25
rect 423 17 425 25
rect 430 17 432 25
rect 440 19 442 25
rect 463 17 465 26
rect 473 17 475 25
rect 480 17 482 25
rect 490 17 492 25
rect 497 17 499 25
rect 507 19 509 25
rect 529 22 531 31
rect 539 25 541 31
rect 549 25 551 31
rect 572 14 574 26
rect 579 14 581 26
rect 589 17 591 26
rect 599 17 601 26
rect 615 22 617 31
<< pmos >>
rect 13 43 15 61
rect 26 50 28 71
rect 33 50 35 71
rect 62 44 64 62
rect 72 51 74 64
rect 82 51 84 64
rect 110 44 112 71
rect 126 44 128 62
rect 136 44 138 62
rect 146 44 148 71
rect 176 44 178 62
rect 186 51 188 64
rect 196 51 198 64
rect 224 44 226 71
rect 240 44 242 62
rect 250 44 252 62
rect 260 44 262 71
rect 287 51 289 64
rect 297 51 299 64
rect 307 44 309 62
rect 339 55 341 71
rect 346 55 348 71
rect 356 55 358 71
rect 363 55 365 71
rect 329 43 331 51
rect 373 53 375 71
rect 396 53 398 71
rect 406 55 408 71
rect 413 55 415 71
rect 423 55 425 71
rect 430 55 432 71
rect 463 53 465 71
rect 473 55 475 71
rect 480 55 482 71
rect 490 55 492 71
rect 497 55 499 71
rect 440 43 442 51
rect 507 43 509 51
rect 529 43 531 61
rect 542 50 544 71
rect 549 50 551 71
rect 571 44 573 71
rect 581 44 583 62
rect 591 44 593 62
rect 607 44 609 71
<< polyct0 >>
rect 15 36 17 38
rect 64 36 66 38
rect 134 36 136 38
rect 144 37 146 39
rect 178 36 180 38
rect 248 36 250 38
rect 258 37 260 39
rect 305 36 307 38
rect 347 46 349 48
rect 354 30 356 32
rect 422 46 424 48
rect 372 31 374 33
rect 397 31 399 33
rect 415 30 417 32
rect 489 46 491 48
rect 464 31 466 33
rect 482 30 484 32
rect 531 36 533 38
rect 573 37 575 39
rect 583 36 585 38
<< polyct1 >>
rect 35 43 37 45
rect 25 36 27 38
rect 84 44 86 46
rect 97 44 99 46
rect 74 36 76 38
rect 198 44 200 46
rect 211 44 213 46
rect 285 44 287 46
rect 113 31 115 33
rect 188 36 190 38
rect 227 31 229 33
rect 324 56 326 58
rect 295 36 297 38
rect 445 56 447 58
rect 337 36 339 38
rect 364 41 366 43
rect 405 41 407 43
rect 512 56 514 58
rect 432 36 434 38
rect 472 41 474 43
rect 499 36 501 38
rect 551 43 553 45
rect 620 44 622 46
rect 541 36 543 38
rect 604 31 606 33
<< ndifct0 >>
rect 28 27 30 29
rect 19 14 21 16
rect 97 27 99 29
rect 87 20 89 22
rect 111 19 113 21
rect 38 14 40 16
rect 123 22 125 24
rect 211 27 213 29
rect 201 20 203 22
rect 225 19 227 21
rect 237 22 239 24
rect 282 20 284 22
rect 324 21 326 23
rect 334 21 336 23
rect 351 19 353 21
rect 368 19 370 21
rect 401 19 403 21
rect 418 19 420 21
rect 435 21 437 23
rect 445 21 447 23
rect 468 19 470 21
rect 485 19 487 21
rect 502 21 504 23
rect 512 21 514 23
rect 544 27 546 29
rect 535 14 537 16
rect 554 14 556 16
rect 594 22 596 24
rect 620 27 622 29
rect 606 19 608 21
<< ndifct1 >>
rect 8 27 10 29
rect 57 22 59 24
rect 133 20 135 22
rect 68 10 70 12
rect 171 22 173 24
rect 151 10 153 12
rect 247 20 249 22
rect 182 10 184 12
rect 312 22 314 24
rect 265 10 267 12
rect 301 10 303 12
rect 378 22 380 24
rect 391 22 393 24
rect 458 22 460 24
rect 524 27 526 29
rect 584 20 586 22
rect 566 10 568 12
<< ntiect1 >>
rect 9 70 11 72
rect 58 70 60 72
rect 131 70 133 72
rect 172 70 174 72
rect 245 70 247 72
rect 311 70 313 72
rect 525 70 527 72
rect 586 70 588 72
<< ptiect1 >>
rect 9 10 11 12
rect 58 10 60 12
rect 98 10 100 12
rect 172 10 174 12
rect 212 10 214 12
rect 311 10 313 12
rect 525 10 527 12
rect 619 10 621 12
<< pdifct0 >>
rect 19 67 21 69
rect 38 60 40 62
rect 67 58 69 60
rect 77 60 79 62
rect 77 53 79 55
rect 87 60 89 62
rect 105 46 107 48
rect 115 67 117 69
rect 115 60 117 62
rect 131 53 133 55
rect 131 46 133 48
rect 151 61 153 63
rect 181 58 183 60
rect 191 60 193 62
rect 191 53 193 55
rect 201 60 203 62
rect 219 46 221 48
rect 229 67 231 69
rect 229 60 231 62
rect 245 53 247 55
rect 245 46 247 48
rect 334 67 336 69
rect 265 61 267 63
rect 282 60 284 62
rect 292 60 294 62
rect 292 53 294 55
rect 302 58 304 60
rect 351 57 353 59
rect 368 67 370 69
rect 324 45 326 47
rect 401 67 403 69
rect 418 57 420 59
rect 435 67 437 69
rect 468 67 470 69
rect 485 57 487 59
rect 502 67 504 69
rect 535 67 537 69
rect 445 45 447 47
rect 512 45 514 47
rect 554 60 556 62
rect 566 61 568 63
rect 602 67 604 69
rect 586 53 588 55
rect 586 46 588 48
rect 602 60 604 62
rect 612 46 614 48
<< pdifct1 >>
rect 8 57 10 59
rect 8 50 10 52
rect 57 53 59 55
rect 57 46 59 48
rect 141 53 143 55
rect 171 53 173 55
rect 171 46 173 48
rect 255 53 257 55
rect 312 53 314 55
rect 312 46 314 48
rect 378 60 380 62
rect 391 60 393 62
rect 458 60 460 62
rect 524 57 526 59
rect 524 50 526 52
rect 576 53 578 55
<< alu0 >>
rect 17 67 19 69
rect 21 67 23 69
rect 17 66 23 67
rect 25 62 42 63
rect 25 60 38 62
rect 40 60 42 62
rect 25 59 42 60
rect 65 60 71 69
rect 10 48 11 59
rect 25 55 29 59
rect 65 58 67 60
rect 69 58 71 60
rect 65 57 71 58
rect 76 62 80 64
rect 76 60 77 62
rect 79 60 80 62
rect 14 51 29 55
rect 76 55 80 60
rect 85 62 91 69
rect 114 67 115 69
rect 117 67 118 69
rect 85 60 87 62
rect 89 60 91 62
rect 85 59 91 60
rect 114 62 118 67
rect 114 60 115 62
rect 117 60 118 62
rect 114 58 118 60
rect 122 63 155 64
rect 122 61 151 63
rect 153 61 155 63
rect 122 60 155 61
rect 179 60 185 69
rect 76 54 77 55
rect 14 38 18 51
rect 63 53 77 54
rect 79 53 80 55
rect 63 50 80 53
rect 33 42 39 43
rect 14 36 15 38
rect 17 36 18 38
rect 14 30 18 36
rect 14 29 32 30
rect 14 27 28 29
rect 30 27 32 29
rect 14 26 32 27
rect 63 38 67 50
rect 122 49 126 60
rect 179 58 181 60
rect 183 58 185 60
rect 179 57 185 58
rect 190 62 194 64
rect 190 60 191 62
rect 193 60 194 62
rect 103 48 126 49
rect 103 46 105 48
rect 107 46 126 48
rect 103 45 126 46
rect 103 39 107 45
rect 63 36 64 38
rect 66 36 67 38
rect 63 31 67 36
rect 63 27 75 31
rect 59 24 60 26
rect 71 23 75 27
rect 96 35 107 39
rect 96 29 100 35
rect 122 39 126 45
rect 130 55 134 57
rect 130 53 131 55
rect 133 53 134 55
rect 130 48 134 53
rect 130 46 131 48
rect 133 47 134 48
rect 133 46 146 47
rect 130 43 146 46
rect 142 41 146 43
rect 142 39 147 41
rect 122 38 138 39
rect 122 36 134 38
rect 136 36 138 38
rect 122 35 138 36
rect 142 37 144 39
rect 146 37 147 39
rect 142 35 147 37
rect 96 27 97 29
rect 99 27 100 29
rect 96 25 100 27
rect 142 31 146 35
rect 122 27 146 31
rect 122 24 126 27
rect 71 22 91 23
rect 122 22 123 24
rect 125 22 126 24
rect 71 20 87 22
rect 89 20 91 22
rect 71 19 91 20
rect 109 21 115 22
rect 109 19 111 21
rect 113 19 115 21
rect 122 20 126 22
rect 190 55 194 60
rect 199 62 205 69
rect 228 67 229 69
rect 231 67 232 69
rect 199 60 201 62
rect 203 60 205 62
rect 199 59 205 60
rect 228 62 232 67
rect 228 60 229 62
rect 231 60 232 62
rect 228 58 232 60
rect 236 63 269 64
rect 236 61 265 63
rect 267 61 269 63
rect 236 60 269 61
rect 280 62 286 69
rect 280 60 282 62
rect 284 60 286 62
rect 190 54 191 55
rect 177 53 191 54
rect 193 53 194 55
rect 177 50 194 53
rect 177 38 181 50
rect 236 49 240 60
rect 280 59 286 60
rect 291 62 295 64
rect 291 60 292 62
rect 294 60 295 62
rect 217 48 240 49
rect 217 46 219 48
rect 221 46 240 48
rect 217 45 240 46
rect 217 39 221 45
rect 177 36 178 38
rect 180 36 181 38
rect 177 31 181 36
rect 177 27 189 31
rect 173 24 174 26
rect 17 16 23 17
rect 17 14 19 16
rect 21 14 23 16
rect 17 13 23 14
rect 36 16 42 17
rect 36 14 38 16
rect 40 14 42 16
rect 36 13 42 14
rect 109 13 115 19
rect 185 23 189 27
rect 210 35 221 39
rect 210 29 214 35
rect 236 39 240 45
rect 244 55 248 57
rect 244 53 245 55
rect 247 53 248 55
rect 244 48 248 53
rect 244 46 245 48
rect 247 47 248 48
rect 247 46 260 47
rect 244 43 260 46
rect 256 41 260 43
rect 291 55 295 60
rect 300 60 306 69
rect 333 67 334 69
rect 336 67 337 69
rect 333 65 337 67
rect 366 67 368 69
rect 370 67 372 69
rect 366 66 372 67
rect 399 67 401 69
rect 403 67 405 69
rect 399 66 405 67
rect 434 67 435 69
rect 437 67 438 69
rect 434 65 438 67
rect 466 67 468 69
rect 470 67 472 69
rect 466 66 472 67
rect 501 67 502 69
rect 504 67 505 69
rect 501 65 505 67
rect 533 67 535 69
rect 537 67 539 69
rect 533 66 539 67
rect 601 67 602 69
rect 604 67 605 69
rect 300 58 302 60
rect 304 58 306 60
rect 300 57 306 58
rect 291 53 292 55
rect 294 54 295 55
rect 294 53 308 54
rect 291 50 308 53
rect 256 39 261 41
rect 236 38 252 39
rect 236 36 248 38
rect 250 36 252 38
rect 236 35 252 36
rect 256 37 258 39
rect 260 37 261 39
rect 256 35 261 37
rect 210 27 211 29
rect 213 27 214 29
rect 210 25 214 27
rect 256 31 260 35
rect 236 27 260 31
rect 236 24 240 27
rect 185 22 205 23
rect 236 22 237 24
rect 239 22 240 24
rect 304 38 308 50
rect 349 59 362 60
rect 349 57 351 59
rect 353 57 362 59
rect 349 56 362 57
rect 358 52 374 56
rect 346 48 350 50
rect 304 36 305 38
rect 307 36 308 38
rect 304 31 308 36
rect 296 27 308 31
rect 296 23 300 27
rect 311 24 312 26
rect 185 20 201 22
rect 203 20 205 22
rect 185 19 205 20
rect 223 21 229 22
rect 223 19 225 21
rect 227 19 229 21
rect 236 20 240 22
rect 280 22 300 23
rect 280 20 282 22
rect 284 20 300 22
rect 280 19 300 20
rect 223 13 229 19
rect 322 47 347 48
rect 322 45 324 47
rect 326 46 347 47
rect 349 46 350 48
rect 326 45 350 46
rect 322 44 350 45
rect 322 24 326 44
rect 346 34 350 44
rect 366 39 367 45
rect 370 35 374 52
rect 346 32 357 34
rect 346 30 354 32
rect 356 30 357 32
rect 370 33 375 35
rect 370 31 372 33
rect 374 31 375 33
rect 346 28 357 30
rect 360 29 375 31
rect 360 27 374 29
rect 322 23 328 24
rect 322 21 324 23
rect 326 21 328 23
rect 322 20 328 21
rect 332 23 338 24
rect 332 21 334 23
rect 336 21 338 23
rect 360 22 364 27
rect 332 13 338 21
rect 349 21 364 22
rect 349 19 351 21
rect 353 19 364 21
rect 349 18 364 19
rect 367 21 371 23
rect 367 19 368 21
rect 370 19 371 21
rect 367 13 371 19
rect 409 59 422 60
rect 409 57 418 59
rect 420 57 422 59
rect 409 56 422 57
rect 397 52 413 56
rect 397 35 401 52
rect 476 59 489 60
rect 421 48 425 50
rect 404 39 405 45
rect 421 46 422 48
rect 424 47 449 48
rect 424 46 445 47
rect 421 45 445 46
rect 447 45 449 47
rect 421 44 449 45
rect 396 33 401 35
rect 421 34 425 44
rect 396 31 397 33
rect 399 31 401 33
rect 414 32 425 34
rect 396 29 411 31
rect 397 27 411 29
rect 414 30 415 32
rect 417 30 425 32
rect 414 28 425 30
rect 400 21 404 23
rect 400 19 401 21
rect 403 19 404 21
rect 400 13 404 19
rect 407 22 411 27
rect 445 24 449 44
rect 433 23 439 24
rect 407 21 422 22
rect 407 19 418 21
rect 420 19 422 21
rect 407 18 422 19
rect 433 21 435 23
rect 437 21 439 23
rect 433 13 439 21
rect 443 23 449 24
rect 443 21 445 23
rect 447 21 449 23
rect 443 20 449 21
rect 476 57 485 59
rect 487 57 489 59
rect 476 56 489 57
rect 464 52 480 56
rect 464 35 468 52
rect 564 63 597 64
rect 541 62 558 63
rect 541 60 554 62
rect 556 60 558 62
rect 564 61 566 63
rect 568 61 597 63
rect 564 60 597 61
rect 541 59 558 60
rect 488 48 492 50
rect 471 39 472 45
rect 488 46 489 48
rect 491 47 516 48
rect 491 46 512 47
rect 488 45 512 46
rect 514 45 516 47
rect 488 44 516 45
rect 463 33 468 35
rect 488 34 492 44
rect 463 31 464 33
rect 466 31 468 33
rect 481 32 492 34
rect 463 29 478 31
rect 464 27 478 29
rect 481 30 482 32
rect 484 30 492 32
rect 481 28 492 30
rect 467 21 471 23
rect 467 19 468 21
rect 470 19 471 21
rect 467 13 471 19
rect 474 22 478 27
rect 512 24 516 44
rect 526 48 527 59
rect 541 55 545 59
rect 530 51 545 55
rect 530 38 534 51
rect 585 55 589 57
rect 585 53 586 55
rect 588 53 589 55
rect 549 42 555 43
rect 530 36 531 38
rect 533 36 534 38
rect 530 30 534 36
rect 530 29 548 30
rect 530 27 544 29
rect 546 27 548 29
rect 530 26 548 27
rect 585 48 589 53
rect 585 47 586 48
rect 573 46 586 47
rect 588 46 589 48
rect 573 43 589 46
rect 593 49 597 60
rect 601 62 605 67
rect 601 60 602 62
rect 604 60 605 62
rect 601 58 605 60
rect 593 48 616 49
rect 593 46 612 48
rect 614 46 616 48
rect 593 45 616 46
rect 573 41 577 43
rect 572 39 577 41
rect 593 39 597 45
rect 572 37 573 39
rect 575 37 577 39
rect 572 35 577 37
rect 581 38 597 39
rect 581 36 583 38
rect 585 36 597 38
rect 581 35 597 36
rect 500 23 506 24
rect 474 21 489 22
rect 474 19 485 21
rect 487 19 489 21
rect 474 18 489 19
rect 500 21 502 23
rect 504 21 506 23
rect 500 13 506 21
rect 510 23 516 24
rect 510 21 512 23
rect 514 21 516 23
rect 510 20 516 21
rect 573 31 577 35
rect 612 39 616 45
rect 612 35 623 39
rect 573 27 597 31
rect 593 24 597 27
rect 619 29 623 35
rect 619 27 620 29
rect 622 27 623 29
rect 619 25 623 27
rect 593 22 594 24
rect 596 22 597 24
rect 593 20 597 22
rect 604 21 610 22
rect 604 19 606 21
rect 608 19 610 21
rect 533 16 539 17
rect 533 14 535 16
rect 537 14 539 16
rect 533 13 539 14
rect 552 16 558 17
rect 552 14 554 16
rect 556 14 558 16
rect 552 13 558 14
rect 604 13 610 19
<< via1 >>
rect 88 51 90 53
rect 39 36 41 38
rect 97 51 99 53
rect 80 27 82 29
rect 105 27 107 29
rect 152 28 154 30
rect 202 51 204 53
rect 170 36 172 38
rect 211 51 213 53
rect 194 27 196 29
rect 266 43 268 45
rect 219 27 221 29
rect 332 52 334 54
rect 313 28 315 30
rect 330 28 332 30
rect 355 44 357 46
rect 379 36 381 38
rect 406 36 408 38
rect 437 28 439 30
rect 504 52 506 54
rect 480 43 482 45
rect 457 28 459 30
rect 505 28 507 30
rect 523 44 525 46
rect 565 28 567 30
<< labels >>
rlabel alu1 125 9 125 9 6 vss
rlabel alu1 125 73 125 73 6 vdd
rlabel alu1 73 73 73 73 6 vdd
rlabel alu1 73 9 73 9 6 vss
rlabel alu1 239 9 239 9 6 vss
rlabel alu1 239 73 239 73 6 vdd
rlabel alu1 267 33 267 33 1 sum
rlabel alu1 187 73 187 73 6 vdd
rlabel alu1 187 9 187 9 6 vss
rlabel alu1 24 9 24 9 6 vss
rlabel alu1 24 73 24 73 6 vdd
rlabel alu1 73 36 73 36 1 a
rlabel via1 88 51 88 51 1 b
rlabel via1 204 52 204 52 1 cin
rlabel alu1 8 39 8 39 1 cout
rlabel alu1 298 9 298 9 4 vss
rlabel alu1 298 37 298 37 4 a
rlabel alu1 290 33 290 33 4 a
rlabel alu1 290 45 290 45 4 b
rlabel alu1 298 73 298 73 4 vdd
rlabel alu1 282 53 282 53 4 b
rlabel alu1 391 37 391 37 6 z
rlabel alu1 399 61 399 61 6 z
rlabel alu1 419 9 419 9 6 vss
rlabel alu1 419 73 419 73 6 vdd
rlabel via1 356 45 356 45 4 a0
rlabel alu1 364 41 364 41 4 a0
rlabel alu1 352 9 352 9 4 vss
rlabel alu1 340 37 340 37 4 a1
rlabel alu1 352 73 352 73 4 vdd
rlabel alu1 332 29 332 29 4 a1
rlabel alu1 486 9 486 9 6 vss
rlabel alu1 486 73 486 73 6 vdd
rlabel alu1 478 44 478 44 1 a2
rlabel alu1 474 39 474 39 1 a2
rlabel alu1 497 37 497 37 1 a3
rlabel alu1 502 28 502 28 1 a3
rlabel via1 506 53 506 53 1 s1
rlabel alu1 514 61 514 61 1 s1
rlabel via1 332 53 332 53 1 s1
rlabel alu1 324 61 324 61 1 s1
rlabel alu1 447 61 447 61 1 s0
rlabel alu1 540 9 540 9 6 vss
rlabel alu1 540 73 540 73 6 vdd
rlabel alu1 556 53 556 53 6 b
rlabel alu1 556 29 556 29 6 a
rlabel alu1 540 45 540 45 6 b
rlabel alu1 548 45 548 45 6 b
rlabel alu1 548 37 548 37 6 a
rlabel alu1 540 37 540 37 6 a
rlabel alu1 614 29 614 29 4 a
rlabel alu1 622 53 622 53 4 b
rlabel alu1 614 61 614 61 4 b
rlabel alu1 606 33 606 33 4 a
rlabel alu1 594 9 594 9 4 vss
rlabel alu1 594 73 594 73 4 vdd
<< end >>
