magic
tech scmos
timestamp 1607699233
<< ab >>
rect -63 5 0 77
rect 4 5 68 77
rect 72 5 135 77
<< nwell >>
rect -67 37 140 82
<< pwell >>
rect -67 0 140 37
<< poly >>
rect -44 71 -42 75
rect -37 71 -35 75
rect -27 71 -25 75
rect -20 71 -18 75
rect -10 71 -8 75
rect 13 71 15 75
rect 23 71 25 75
rect 30 71 32 75
rect 40 71 42 75
rect 47 71 49 75
rect 80 71 82 75
rect 90 71 92 75
rect 97 71 99 75
rect 107 71 109 75
rect 114 71 116 75
rect -61 58 -55 60
rect -61 56 -59 58
rect -57 56 -55 58
rect -61 54 -52 56
rect -54 51 -52 54
rect -54 25 -52 43
rect -44 40 -42 55
rect -37 50 -35 55
rect -38 48 -32 50
rect -38 46 -36 48
rect -34 46 -32 48
rect -38 44 -32 46
rect -27 40 -25 55
rect -20 45 -18 55
rect 60 58 66 60
rect 60 56 62 58
rect 64 56 66 58
rect -48 38 -42 40
rect -48 36 -46 38
rect -44 36 -42 38
rect -48 34 -42 36
rect -44 25 -42 34
rect -37 38 -25 40
rect -21 43 -15 45
rect -21 41 -19 43
rect -17 41 -15 43
rect -21 39 -15 41
rect -37 25 -35 38
rect -31 32 -25 34
rect -31 30 -29 32
rect -27 30 -25 32
rect -31 28 -25 30
rect -27 25 -25 28
rect -20 25 -18 39
rect -10 35 -8 53
rect 13 35 15 53
rect 23 45 25 55
rect 20 43 26 45
rect 20 41 22 43
rect 24 41 26 43
rect 20 39 26 41
rect 30 40 32 55
rect 40 50 42 55
rect 37 48 43 50
rect 37 46 39 48
rect 41 46 43 48
rect 37 44 43 46
rect 47 40 49 55
rect 57 54 66 56
rect 57 51 59 54
rect 127 58 133 60
rect 127 56 129 58
rect 131 56 133 58
rect -13 33 -7 35
rect -13 31 -11 33
rect -9 31 -7 33
rect -13 29 -7 31
rect 12 33 18 35
rect 12 31 14 33
rect 16 31 18 33
rect 12 29 18 31
rect -10 26 -8 29
rect 13 26 15 29
rect -54 9 -52 19
rect 23 25 25 39
rect 30 38 42 40
rect 30 32 36 34
rect 30 30 32 32
rect 34 30 36 32
rect 30 28 36 30
rect 30 25 32 28
rect 40 25 42 38
rect 47 38 53 40
rect 47 36 49 38
rect 51 36 53 38
rect 47 34 53 36
rect 47 25 49 34
rect 57 25 59 43
rect 80 35 82 53
rect 90 45 92 55
rect 87 43 93 45
rect 87 41 89 43
rect 91 41 93 43
rect 87 39 93 41
rect 97 40 99 55
rect 107 50 109 55
rect 104 48 110 50
rect 104 46 106 48
rect 108 46 110 48
rect 104 44 110 46
rect 114 40 116 55
rect 124 54 133 56
rect 124 51 126 54
rect 79 33 85 35
rect 79 31 81 33
rect 83 31 85 33
rect 79 29 85 31
rect 80 26 82 29
rect -44 13 -42 17
rect -37 9 -35 17
rect -27 12 -25 17
rect -20 12 -18 17
rect -10 12 -8 17
rect 13 12 15 17
rect 23 12 25 17
rect 30 12 32 17
rect -54 7 -35 9
rect 40 9 42 17
rect 47 13 49 17
rect 57 9 59 19
rect 90 25 92 39
rect 97 38 109 40
rect 97 32 103 34
rect 97 30 99 32
rect 101 30 103 32
rect 97 28 103 30
rect 97 25 99 28
rect 107 25 109 38
rect 114 38 120 40
rect 114 36 116 38
rect 118 36 120 38
rect 114 34 120 36
rect 114 25 116 34
rect 124 25 126 43
rect 80 12 82 17
rect 90 12 92 17
rect 97 12 99 17
rect 40 7 59 9
rect 107 9 109 17
rect 114 13 116 17
rect 124 9 126 19
rect 107 7 126 9
<< ndif >>
rect -15 25 -10 26
rect -61 23 -54 25
rect -61 21 -59 23
rect -57 21 -54 23
rect -61 19 -54 21
rect -52 23 -44 25
rect -52 21 -49 23
rect -47 21 -44 23
rect -52 19 -44 21
rect -50 17 -44 19
rect -42 17 -37 25
rect -35 21 -27 25
rect -35 19 -32 21
rect -30 19 -27 21
rect -35 17 -27 19
rect -25 17 -20 25
rect -18 21 -10 25
rect -18 19 -15 21
rect -13 19 -10 21
rect -18 17 -10 19
rect -8 24 -1 26
rect -8 22 -5 24
rect -3 22 -1 24
rect -8 20 -1 22
rect 6 24 13 26
rect 6 22 8 24
rect 10 22 13 24
rect 6 20 13 22
rect -8 17 -3 20
rect 8 17 13 20
rect 15 25 20 26
rect 15 21 23 25
rect 15 19 18 21
rect 20 19 23 21
rect 15 17 23 19
rect 25 17 30 25
rect 32 21 40 25
rect 32 19 35 21
rect 37 19 40 21
rect 32 17 40 19
rect 42 17 47 25
rect 49 23 57 25
rect 49 21 52 23
rect 54 21 57 23
rect 49 19 57 21
rect 59 23 66 25
rect 59 21 62 23
rect 64 21 66 23
rect 59 19 66 21
rect 73 24 80 26
rect 73 22 75 24
rect 77 22 80 24
rect 73 20 80 22
rect 49 17 55 19
rect 75 17 80 20
rect 82 25 87 26
rect 82 21 90 25
rect 82 19 85 21
rect 87 19 90 21
rect 82 17 90 19
rect 92 17 97 25
rect 99 21 107 25
rect 99 19 102 21
rect 104 19 107 21
rect 99 17 107 19
rect 109 17 114 25
rect 116 23 124 25
rect 116 21 119 23
rect 121 21 124 23
rect 116 19 124 21
rect 126 23 133 25
rect 126 21 129 23
rect 131 21 133 23
rect 126 19 133 21
rect 116 17 122 19
<< pdif >>
rect -51 69 -44 71
rect -51 67 -49 69
rect -47 67 -44 69
rect -51 59 -44 67
rect -50 55 -44 59
rect -42 55 -37 71
rect -35 59 -27 71
rect -35 57 -32 59
rect -30 57 -27 59
rect -35 55 -27 57
rect -25 55 -20 71
rect -18 69 -10 71
rect -18 67 -15 69
rect -13 67 -10 69
rect -18 55 -10 67
rect -50 51 -46 55
rect -59 49 -54 51
rect -61 47 -54 49
rect -61 45 -59 47
rect -57 45 -54 47
rect -61 43 -54 45
rect -52 43 -46 51
rect -15 53 -10 55
rect -8 64 -3 71
rect 8 64 13 71
rect -8 62 -1 64
rect -8 60 -5 62
rect -3 60 -1 62
rect -8 58 -1 60
rect 6 62 13 64
rect 6 60 8 62
rect 10 60 13 62
rect 6 58 13 60
rect -8 53 -3 58
rect 8 53 13 58
rect 15 69 23 71
rect 15 67 18 69
rect 20 67 23 69
rect 15 55 23 67
rect 25 55 30 71
rect 32 59 40 71
rect 32 57 35 59
rect 37 57 40 59
rect 32 55 40 57
rect 42 55 47 71
rect 49 69 56 71
rect 49 67 52 69
rect 54 67 56 69
rect 49 59 56 67
rect 75 64 80 71
rect 73 62 80 64
rect 73 60 75 62
rect 77 60 80 62
rect 49 55 55 59
rect 73 58 80 60
rect 15 53 20 55
rect 51 51 55 55
rect 75 53 80 58
rect 82 69 90 71
rect 82 67 85 69
rect 87 67 90 69
rect 82 55 90 67
rect 92 55 97 71
rect 99 59 107 71
rect 99 57 102 59
rect 104 57 107 59
rect 99 55 107 57
rect 109 55 114 71
rect 116 69 123 71
rect 116 67 119 69
rect 121 67 123 69
rect 116 59 123 67
rect 116 55 122 59
rect 82 53 87 55
rect 51 43 57 51
rect 59 49 64 51
rect 59 47 66 49
rect 59 45 62 47
rect 64 45 66 47
rect 59 43 66 45
rect 118 51 122 55
rect 118 43 124 51
rect 126 49 131 51
rect 126 47 133 49
rect 126 45 129 47
rect 131 45 133 47
rect 126 43 133 45
<< alu1 >>
rect -65 69 137 77
rect -61 58 -56 64
rect -14 62 -1 63
rect -14 60 -5 62
rect -3 60 -1 62
rect -61 56 -59 58
rect -57 56 -56 58
rect -14 59 -1 60
rect -61 55 -56 56
rect -61 54 -48 55
rect -61 52 -51 54
rect -49 52 -48 54
rect -61 51 -48 52
rect -47 38 -41 40
rect -47 36 -46 38
rect -44 36 -41 38
rect -47 31 -41 36
rect -54 27 -41 31
rect -29 43 -17 48
rect -29 42 -19 43
rect -21 41 -19 42
rect -21 34 -17 41
rect -5 38 -1 59
rect -5 36 -4 38
rect -2 36 -1 38
rect -5 26 -1 36
rect -6 24 -1 26
rect -6 22 -5 24
rect -3 22 -1 24
rect -6 20 -1 22
rect -5 18 -1 20
rect 6 62 19 63
rect 6 60 8 62
rect 10 60 19 62
rect 6 59 19 60
rect 6 26 10 59
rect 61 58 66 64
rect 61 56 62 58
rect 64 56 66 58
rect 61 55 66 56
rect 53 51 66 55
rect 73 62 86 63
rect 73 60 75 62
rect 77 60 86 62
rect 73 59 86 60
rect 22 43 34 48
rect 24 42 34 43
rect 24 41 26 42
rect 22 38 26 41
rect 22 36 23 38
rect 25 36 26 38
rect 22 34 26 36
rect 46 38 52 40
rect 46 36 49 38
rect 51 36 52 38
rect 46 31 52 36
rect 46 30 59 31
rect 46 28 54 30
rect 56 28 59 30
rect 46 27 59 28
rect 6 24 11 26
rect 6 22 8 24
rect 10 22 11 24
rect 6 20 11 22
rect 6 18 10 20
rect 73 30 77 59
rect 128 58 133 64
rect 128 56 129 58
rect 131 56 133 58
rect 128 55 133 56
rect 120 54 133 55
rect 120 52 121 54
rect 123 52 133 54
rect 120 51 133 52
rect 89 43 101 48
rect 91 42 101 43
rect 91 41 93 42
rect 73 28 74 30
rect 76 28 77 30
rect 89 34 93 41
rect 73 26 77 28
rect 113 38 119 40
rect 113 36 116 38
rect 118 36 119 38
rect 113 31 119 36
rect 113 27 126 31
rect 73 24 78 26
rect 73 22 75 24
rect 77 22 78 24
rect 73 20 78 22
rect 73 18 77 20
rect -65 5 137 13
<< alu2 >>
rect -52 54 125 55
rect -52 52 -51 54
rect -49 52 121 54
rect 123 52 125 54
rect -52 51 125 52
rect -5 38 26 39
rect -5 36 -4 38
rect -2 36 23 38
rect 25 36 26 38
rect -5 35 26 36
rect 53 30 77 31
rect 53 28 54 30
rect 56 28 74 30
rect 76 28 77 30
rect 53 27 77 28
<< nmos >>
rect -54 19 -52 25
rect -44 17 -42 25
rect -37 17 -35 25
rect -27 17 -25 25
rect -20 17 -18 25
rect -10 17 -8 26
rect 13 17 15 26
rect 23 17 25 25
rect 30 17 32 25
rect 40 17 42 25
rect 47 17 49 25
rect 57 19 59 25
rect 80 17 82 26
rect 90 17 92 25
rect 97 17 99 25
rect 107 17 109 25
rect 114 17 116 25
rect 124 19 126 25
<< pmos >>
rect -44 55 -42 71
rect -37 55 -35 71
rect -27 55 -25 71
rect -20 55 -18 71
rect -54 43 -52 51
rect -10 53 -8 71
rect 13 53 15 71
rect 23 55 25 71
rect 30 55 32 71
rect 40 55 42 71
rect 47 55 49 71
rect 80 53 82 71
rect 90 55 92 71
rect 97 55 99 71
rect 107 55 109 71
rect 114 55 116 71
rect 57 43 59 51
rect 124 43 126 51
<< polyct0 >>
rect -36 46 -34 48
rect -29 30 -27 32
rect 39 46 41 48
rect -11 31 -9 33
rect 14 31 16 33
rect 32 30 34 32
rect 106 46 108 48
rect 81 31 83 33
rect 99 30 101 32
<< polyct1 >>
rect -59 56 -57 58
rect 62 56 64 58
rect -46 36 -44 38
rect -19 41 -17 43
rect 22 41 24 43
rect 129 56 131 58
rect 49 36 51 38
rect 89 41 91 43
rect 116 36 118 38
<< ndifct0 >>
rect -59 21 -57 23
rect -49 21 -47 23
rect -32 19 -30 21
rect -15 19 -13 21
rect 18 19 20 21
rect 35 19 37 21
rect 52 21 54 23
rect 62 21 64 23
rect 85 19 87 21
rect 102 19 104 21
rect 119 21 121 23
rect 129 21 131 23
<< ndifct1 >>
rect -5 22 -3 24
rect 8 22 10 24
rect 75 22 77 24
<< pdifct0 >>
rect -49 67 -47 69
rect -32 57 -30 59
rect -15 67 -13 69
rect -59 45 -57 47
rect 18 67 20 69
rect 35 57 37 59
rect 52 67 54 69
rect 85 67 87 69
rect 102 57 104 59
rect 119 67 121 69
rect 62 45 64 47
rect 129 45 131 47
<< pdifct1 >>
rect -5 60 -3 62
rect 8 60 10 62
rect 75 60 77 62
<< alu0 >>
rect -50 67 -49 69
rect -47 67 -46 69
rect -50 65 -46 67
rect -17 67 -15 69
rect -13 67 -11 69
rect -17 66 -11 67
rect 16 67 18 69
rect 20 67 22 69
rect 16 66 22 67
rect 51 67 52 69
rect 54 67 55 69
rect 51 65 55 67
rect 83 67 85 69
rect 87 67 89 69
rect 83 66 89 67
rect 118 67 119 69
rect 121 67 122 69
rect 118 65 122 67
rect -34 59 -21 60
rect -34 57 -32 59
rect -30 57 -21 59
rect -34 56 -21 57
rect -25 52 -9 56
rect -37 48 -33 50
rect -61 47 -36 48
rect -61 45 -59 47
rect -57 46 -36 47
rect -34 46 -33 48
rect -57 45 -33 46
rect -61 44 -33 45
rect -61 24 -57 44
rect -37 34 -33 44
rect -17 39 -16 45
rect -13 35 -9 52
rect -37 32 -26 34
rect -37 30 -29 32
rect -27 30 -26 32
rect -13 33 -8 35
rect -13 31 -11 33
rect -9 31 -8 33
rect -37 28 -26 30
rect -23 29 -8 31
rect -23 27 -9 29
rect -61 23 -55 24
rect -61 21 -59 23
rect -57 21 -55 23
rect -61 20 -55 21
rect -51 23 -45 24
rect -51 21 -49 23
rect -47 21 -45 23
rect -23 22 -19 27
rect -51 13 -45 21
rect -34 21 -19 22
rect -34 19 -32 21
rect -30 19 -19 21
rect -34 18 -19 19
rect -16 21 -12 23
rect -16 19 -15 21
rect -13 19 -12 21
rect -16 13 -12 19
rect 26 59 39 60
rect 26 57 35 59
rect 37 57 39 59
rect 26 56 39 57
rect 14 52 30 56
rect 14 35 18 52
rect 93 59 106 60
rect 38 48 42 50
rect 21 39 22 45
rect 38 46 39 48
rect 41 47 66 48
rect 41 46 62 47
rect 38 45 62 46
rect 64 45 66 47
rect 38 44 66 45
rect 13 33 18 35
rect 38 34 42 44
rect 13 31 14 33
rect 16 31 18 33
rect 31 32 42 34
rect 13 29 28 31
rect 14 27 28 29
rect 31 30 32 32
rect 34 30 42 32
rect 31 28 42 30
rect 17 21 21 23
rect 17 19 18 21
rect 20 19 21 21
rect 17 13 21 19
rect 24 22 28 27
rect 62 24 66 44
rect 50 23 56 24
rect 24 21 39 22
rect 24 19 35 21
rect 37 19 39 21
rect 24 18 39 19
rect 50 21 52 23
rect 54 21 56 23
rect 50 13 56 21
rect 60 23 66 24
rect 60 21 62 23
rect 64 21 66 23
rect 60 20 66 21
rect 93 57 102 59
rect 104 57 106 59
rect 93 56 106 57
rect 81 52 97 56
rect 81 35 85 52
rect 105 48 109 50
rect 88 39 89 45
rect 105 46 106 48
rect 108 47 133 48
rect 108 46 129 47
rect 105 45 129 46
rect 131 45 133 47
rect 105 44 133 45
rect 80 33 85 35
rect 105 34 109 44
rect 80 31 81 33
rect 83 31 85 33
rect 98 32 109 34
rect 80 29 95 31
rect 81 27 95 29
rect 98 30 99 32
rect 101 30 109 32
rect 98 28 109 30
rect 84 21 88 23
rect 84 19 85 21
rect 87 19 88 21
rect 84 13 88 19
rect 91 22 95 27
rect 129 24 133 44
rect 117 23 123 24
rect 91 21 106 22
rect 91 19 102 21
rect 104 19 106 21
rect 91 18 106 19
rect 117 21 119 23
rect 121 21 123 23
rect 117 13 123 21
rect 127 23 133 24
rect 127 21 129 23
rect 131 21 133 23
rect 127 20 133 21
<< via1 >>
rect -51 52 -49 54
rect -4 36 -2 38
rect 23 36 25 38
rect 54 28 56 30
rect 121 52 123 54
rect 74 28 76 30
<< labels >>
rlabel alu1 8 37 8 37 6 z
rlabel alu1 16 61 16 61 6 z
rlabel alu1 36 9 36 9 6 vss
rlabel alu1 36 73 36 73 6 vdd
rlabel alu1 -27 45 -27 45 4 a0
rlabel alu1 -19 41 -19 41 4 a0
rlabel alu1 -31 9 -31 9 4 vss
rlabel alu1 -43 37 -43 37 4 a1
rlabel alu1 -31 73 -31 73 4 vdd
rlabel alu1 -51 29 -51 29 4 a1
rlabel alu0 103 31 103 31 6 sn
rlabel alu1 103 9 103 9 6 vss
rlabel alu1 103 73 103 73 6 vdd
rlabel alu1 95 44 95 44 1 a2
rlabel alu1 91 39 91 39 1 a2
rlabel alu1 114 37 114 37 1 a3
rlabel alu1 119 28 119 28 1 a3
rlabel via1 123 53 123 53 1 s1
rlabel alu1 131 61 131 61 1 s1
rlabel via1 -51 53 -51 53 1 s1
rlabel alu1 -59 61 -59 61 1 s1
rlabel alu1 64 61 64 61 1 s0
<< end >>
