magic
tech scmos
timestamp 1608791518
<< ab >>
rect -35 5 45 77
rect 47 5 150 77
rect 152 5 215 77
<< nwell >>
rect -40 37 220 82
<< pwell >>
rect -40 0 220 37
<< poly >>
rect -13 71 -11 75
rect -6 71 -4 75
rect -26 61 -24 66
rect 63 71 65 75
rect 14 62 16 66
rect 24 64 26 69
rect 34 64 36 69
rect -26 40 -24 43
rect -13 40 -11 50
rect -6 47 -4 50
rect -6 45 0 47
rect -6 43 -4 45
rect -2 43 0 45
rect -6 41 0 43
rect -26 38 -20 40
rect -26 36 -24 38
rect -22 36 -20 38
rect -26 34 -20 36
rect -16 38 -10 40
rect -16 36 -14 38
rect -12 36 -10 38
rect -16 34 -10 36
rect -26 31 -24 34
rect -16 31 -14 34
rect -6 31 -4 41
rect 14 40 16 44
rect 24 40 26 51
rect 34 48 36 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 48 46 54 48
rect 48 44 50 46
rect 52 44 54 46
rect 99 71 101 75
rect 79 62 81 66
rect 89 62 91 66
rect 168 71 170 75
rect 119 62 121 66
rect 129 64 131 69
rect 139 64 141 69
rect 48 42 54 44
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 29 16 34
rect 27 29 29 34
rect 34 29 36 42
rect 52 41 54 42
rect 63 41 65 44
rect 79 41 81 44
rect 52 39 65 41
rect 71 39 81 41
rect 89 40 91 44
rect 99 41 101 44
rect 55 31 57 39
rect 71 35 73 39
rect 64 33 73 35
rect 85 38 91 40
rect 85 36 87 38
rect 89 36 91 38
rect 85 34 91 36
rect 95 39 101 41
rect 95 37 97 39
rect 99 37 101 39
rect 95 35 101 37
rect 119 40 121 44
rect 129 40 131 51
rect 139 48 141 51
rect 139 46 145 48
rect 139 44 141 46
rect 143 44 145 46
rect 139 42 145 44
rect 153 46 159 48
rect 153 44 155 46
rect 157 44 159 46
rect 204 71 206 75
rect 184 62 186 66
rect 194 62 196 66
rect 153 42 159 44
rect 119 38 125 40
rect 119 36 121 38
rect 123 36 125 38
rect 64 31 66 33
rect 68 31 73 33
rect -26 17 -24 22
rect -16 20 -14 25
rect -6 20 -4 25
rect 14 16 16 20
rect 64 29 73 31
rect 89 31 91 34
rect 71 26 73 29
rect 81 26 83 30
rect 89 29 93 31
rect 91 26 93 29
rect 98 26 100 35
rect 119 34 125 36
rect 129 38 135 40
rect 129 36 131 38
rect 133 36 135 38
rect 129 34 135 36
rect 119 29 121 34
rect 132 29 134 34
rect 139 29 141 42
rect 157 41 159 42
rect 168 41 170 44
rect 184 41 186 44
rect 157 39 170 41
rect 176 39 186 41
rect 194 40 196 44
rect 204 41 206 44
rect 160 31 162 39
rect 176 35 178 39
rect 169 33 178 35
rect 190 38 196 40
rect 190 36 192 38
rect 194 36 196 38
rect 190 34 196 36
rect 200 39 206 41
rect 200 37 202 39
rect 204 37 206 39
rect 200 35 206 37
rect 169 31 171 33
rect 173 31 178 33
rect 55 19 57 22
rect 27 13 29 18
rect 34 13 36 18
rect 55 17 60 19
rect 58 9 60 17
rect 71 13 73 17
rect 81 9 83 17
rect 119 16 121 20
rect 169 29 178 31
rect 194 31 196 34
rect 176 26 178 29
rect 186 26 188 30
rect 194 29 198 31
rect 196 26 198 29
rect 203 26 205 35
rect 160 19 162 22
rect 91 9 93 14
rect 98 9 100 14
rect 58 7 83 9
rect 132 13 134 18
rect 139 13 141 18
rect 160 17 165 19
rect 163 9 165 17
rect 176 13 178 17
rect 186 9 188 17
rect 196 9 198 14
rect 203 9 205 14
rect 163 7 188 9
<< ndif >>
rect -33 29 -26 31
rect -33 27 -31 29
rect -29 27 -26 29
rect -33 25 -26 27
rect -31 22 -26 25
rect -24 25 -16 31
rect -14 29 -6 31
rect -14 27 -11 29
rect -9 27 -6 29
rect -14 25 -6 27
rect -4 25 3 31
rect 48 29 55 31
rect 9 26 14 29
rect -24 22 -18 25
rect -22 18 -18 22
rect -2 18 3 25
rect 7 24 14 26
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 20 27 29
rect -22 16 -16 18
rect -22 14 -20 16
rect -18 14 -16 16
rect -22 12 -16 14
rect -3 16 3 18
rect 18 18 27 20
rect 29 18 34 29
rect 36 24 41 29
rect 48 27 50 29
rect 52 27 55 29
rect 48 25 55 27
rect 36 22 43 24
rect 50 22 55 25
rect 57 26 62 31
rect 153 29 160 31
rect 114 26 119 29
rect 57 22 71 26
rect 36 20 39 22
rect 41 20 43 22
rect 36 18 43 20
rect 62 21 71 22
rect 62 19 64 21
rect 66 19 71 21
rect -3 14 -1 16
rect 1 14 3 16
rect -3 12 3 14
rect 18 12 25 18
rect 62 17 71 19
rect 73 24 81 26
rect 73 22 76 24
rect 78 22 81 24
rect 73 17 81 22
rect 83 22 91 26
rect 83 20 86 22
rect 88 20 91 22
rect 83 17 91 20
rect 18 10 20 12
rect 22 10 25 12
rect 18 8 25 10
rect 86 14 91 17
rect 93 14 98 26
rect 100 14 108 26
rect 112 24 119 26
rect 112 22 114 24
rect 116 22 119 24
rect 112 20 119 22
rect 121 20 132 29
rect 123 18 132 20
rect 134 18 139 29
rect 141 24 146 29
rect 153 27 155 29
rect 157 27 160 29
rect 153 25 160 27
rect 141 22 148 24
rect 155 22 160 25
rect 162 26 167 31
rect 162 22 176 26
rect 141 20 144 22
rect 146 20 148 22
rect 141 18 148 20
rect 167 21 176 22
rect 167 19 169 21
rect 171 19 176 21
rect 102 12 108 14
rect 102 10 104 12
rect 106 10 108 12
rect 102 8 108 10
rect 123 12 130 18
rect 167 17 176 19
rect 178 24 186 26
rect 178 22 181 24
rect 183 22 186 24
rect 178 17 186 22
rect 188 22 196 26
rect 188 20 191 22
rect 193 20 196 22
rect 188 17 196 20
rect 123 10 125 12
rect 127 10 130 12
rect 123 8 130 10
rect 191 14 196 17
rect 198 14 203 26
rect 205 14 213 26
rect 207 12 213 14
rect 207 10 209 12
rect 211 10 213 12
rect 207 8 213 10
<< pdif >>
rect -22 69 -13 71
rect -22 67 -20 69
rect -18 67 -13 69
rect -22 61 -13 67
rect -33 59 -26 61
rect -33 57 -31 59
rect -29 57 -26 59
rect -33 52 -26 57
rect -33 50 -31 52
rect -29 50 -26 52
rect -33 48 -26 50
rect -31 43 -26 48
rect -24 50 -13 61
rect -11 50 -6 71
rect -4 64 1 71
rect -4 62 3 64
rect 18 62 24 64
rect -4 60 -1 62
rect 1 60 3 62
rect -4 58 3 60
rect -4 50 1 58
rect 9 57 14 62
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect -24 43 -16 50
rect 7 48 14 53
rect 7 46 9 48
rect 11 46 14 48
rect 7 44 14 46
rect 16 60 24 62
rect 16 58 19 60
rect 21 58 24 60
rect 16 51 24 58
rect 26 62 34 64
rect 26 60 29 62
rect 31 60 34 62
rect 26 55 34 60
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 62 43 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 51 43 60
rect 16 44 22 51
rect 58 50 63 71
rect 56 48 63 50
rect 56 46 58 48
rect 60 46 63 48
rect 56 44 63 46
rect 65 69 77 71
rect 65 67 68 69
rect 70 67 77 69
rect 65 62 77 67
rect 94 62 99 71
rect 65 60 68 62
rect 70 60 79 62
rect 65 44 79 60
rect 81 55 89 62
rect 81 53 84 55
rect 86 53 89 55
rect 81 48 89 53
rect 81 46 84 48
rect 86 46 89 48
rect 81 44 89 46
rect 91 55 99 62
rect 91 53 94 55
rect 96 53 99 55
rect 91 44 99 53
rect 101 65 106 71
rect 101 63 108 65
rect 101 61 104 63
rect 106 61 108 63
rect 123 62 129 64
rect 101 59 108 61
rect 101 44 106 59
rect 114 57 119 62
rect 112 55 119 57
rect 112 53 114 55
rect 116 53 119 55
rect 112 48 119 53
rect 112 46 114 48
rect 116 46 119 48
rect 112 44 119 46
rect 121 60 129 62
rect 121 58 124 60
rect 126 58 129 60
rect 121 51 129 58
rect 131 62 139 64
rect 131 60 134 62
rect 136 60 139 62
rect 131 55 139 60
rect 131 53 134 55
rect 136 53 139 55
rect 131 51 139 53
rect 141 62 148 64
rect 141 60 144 62
rect 146 60 148 62
rect 141 51 148 60
rect 121 44 127 51
rect 163 50 168 71
rect 161 48 168 50
rect 161 46 163 48
rect 165 46 168 48
rect 161 44 168 46
rect 170 69 182 71
rect 170 67 173 69
rect 175 67 182 69
rect 170 62 182 67
rect 199 62 204 71
rect 170 60 173 62
rect 175 60 184 62
rect 170 44 184 60
rect 186 55 194 62
rect 186 53 189 55
rect 191 53 194 55
rect 186 48 194 53
rect 186 46 189 48
rect 191 46 194 48
rect 186 44 194 46
rect 196 55 204 62
rect 196 53 199 55
rect 201 53 204 55
rect 196 44 204 53
rect 206 65 211 71
rect 206 63 213 65
rect 206 61 209 63
rect 211 61 213 63
rect 206 59 213 61
rect 206 44 211 59
<< alu1 >>
rect -37 72 217 77
rect -37 70 -30 72
rect -28 70 10 72
rect 12 70 84 72
rect 86 70 115 72
rect 117 70 189 72
rect 191 70 217 72
rect -37 69 217 70
rect -33 63 -29 64
rect -33 59 -20 63
rect -33 57 -31 59
rect -33 52 -29 57
rect -33 50 -31 52
rect -33 31 -29 50
rect -1 55 3 56
rect -1 53 0 55
rect 2 53 3 55
rect -1 47 3 53
rect -18 45 3 47
rect -18 43 -4 45
rect -2 43 3 45
rect 7 55 12 57
rect 7 53 9 55
rect 11 53 12 55
rect 48 58 60 64
rect 7 48 12 53
rect 7 46 9 48
rect 11 46 12 48
rect 7 44 12 46
rect 7 39 11 44
rect -33 29 -28 31
rect -33 27 -31 29
rect -29 27 -28 29
rect -33 25 -28 27
rect -18 38 11 39
rect -18 36 -14 38
rect -12 36 11 38
rect -18 35 11 36
rect -1 26 3 35
rect 7 24 11 35
rect 39 49 43 56
rect 48 49 53 58
rect 39 47 53 49
rect 30 46 53 47
rect 30 44 36 46
rect 38 44 50 46
rect 52 44 53 46
rect 30 43 43 44
rect 47 43 53 44
rect 48 42 53 43
rect 22 38 36 39
rect 22 36 26 38
rect 28 36 36 38
rect 22 35 36 36
rect 7 22 9 24
rect 11 22 19 24
rect 7 18 19 22
rect 31 29 36 35
rect 31 27 32 29
rect 34 27 36 29
rect 31 26 36 27
rect 64 33 69 40
rect 92 55 108 56
rect 92 53 94 55
rect 96 53 108 55
rect 92 51 108 53
rect 64 32 66 33
rect 56 31 66 32
rect 68 31 69 33
rect 56 29 69 31
rect 56 27 59 29
rect 61 27 69 29
rect 56 26 69 27
rect 104 29 108 51
rect 104 27 105 29
rect 107 27 108 29
rect 104 23 108 27
rect 84 22 108 23
rect 84 20 86 22
rect 88 20 108 22
rect 84 19 108 20
rect 112 55 117 57
rect 112 53 114 55
rect 116 53 117 55
rect 153 58 165 64
rect 112 48 117 53
rect 112 46 114 48
rect 116 46 117 48
rect 112 44 117 46
rect 112 24 116 44
rect 144 49 148 56
rect 153 49 158 58
rect 144 47 158 49
rect 135 46 158 47
rect 135 44 141 46
rect 143 44 155 46
rect 157 44 158 46
rect 135 43 148 44
rect 152 43 158 44
rect 153 42 158 43
rect 127 38 141 39
rect 127 36 131 38
rect 133 36 141 38
rect 127 35 141 36
rect 112 22 114 24
rect 116 22 124 24
rect 112 18 124 22
rect 136 29 141 35
rect 136 27 137 29
rect 139 27 141 29
rect 136 26 141 27
rect 169 33 174 40
rect 197 55 213 56
rect 197 53 199 55
rect 201 53 213 55
rect 197 51 213 53
rect 169 32 171 33
rect 161 31 171 32
rect 173 31 174 33
rect 161 29 174 31
rect 161 27 164 29
rect 166 27 174 29
rect 161 26 174 27
rect 209 23 213 51
rect 189 22 213 23
rect 189 20 191 22
rect 193 20 213 22
rect 189 19 213 20
rect -37 12 217 13
rect -37 10 -30 12
rect -28 10 10 12
rect 12 10 20 12
rect 22 10 51 12
rect 53 10 104 12
rect 106 10 115 12
rect 117 10 125 12
rect 127 10 156 12
rect 158 10 209 12
rect 211 10 217 12
rect -37 5 217 10
<< alu2 >>
rect -1 55 117 56
rect -1 53 0 55
rect 2 53 114 55
rect 116 53 117 55
rect -1 52 117 53
rect 31 29 64 30
rect 31 27 32 29
rect 34 27 59 29
rect 61 27 64 29
rect 31 26 64 27
rect 104 29 169 30
rect 104 27 105 29
rect 107 27 137 29
rect 139 27 164 29
rect 166 27 169 29
rect 104 26 169 27
<< ptie >>
rect -32 12 -26 14
rect 8 12 14 14
rect -32 10 -30 12
rect -28 10 -26 12
rect -32 8 -26 10
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 49 12 55 14
rect 49 10 51 12
rect 53 10 55 12
rect 49 8 55 10
rect 113 12 119 14
rect 113 10 115 12
rect 117 10 119 12
rect 113 8 119 10
rect 154 12 160 14
rect 154 10 156 12
rect 158 10 160 12
rect 154 8 160 10
<< ntie >>
rect -32 72 -26 74
rect -32 70 -30 72
rect -28 70 -26 72
rect 8 72 14 74
rect -32 68 -26 70
rect 8 70 10 72
rect 12 70 14 72
rect 82 72 88 74
rect 8 68 14 70
rect 82 70 84 72
rect 86 70 88 72
rect 113 72 119 74
rect 82 68 88 70
rect 113 70 115 72
rect 117 70 119 72
rect 187 72 193 74
rect 113 68 119 70
rect 187 70 189 72
rect 191 70 193 72
rect 187 68 193 70
<< nmos >>
rect -26 22 -24 31
rect -16 25 -14 31
rect -6 25 -4 31
rect 14 20 16 29
rect 27 18 29 29
rect 34 18 36 29
rect 55 22 57 31
rect 71 17 73 26
rect 81 17 83 26
rect 91 14 93 26
rect 98 14 100 26
rect 119 20 121 29
rect 132 18 134 29
rect 139 18 141 29
rect 160 22 162 31
rect 176 17 178 26
rect 186 17 188 26
rect 196 14 198 26
rect 203 14 205 26
<< pmos >>
rect -26 43 -24 61
rect -13 50 -11 71
rect -6 50 -4 71
rect 14 44 16 62
rect 24 51 26 64
rect 34 51 36 64
rect 63 44 65 71
rect 79 44 81 62
rect 89 44 91 62
rect 99 44 101 71
rect 119 44 121 62
rect 129 51 131 64
rect 139 51 141 64
rect 168 44 170 71
rect 184 44 186 62
rect 194 44 196 62
rect 204 44 206 71
<< polyct0 >>
rect -24 36 -22 38
rect 16 36 18 38
rect 87 36 89 38
rect 97 37 99 39
rect 121 36 123 38
rect 192 36 194 38
rect 202 37 204 39
<< polyct1 >>
rect -4 43 -2 45
rect -14 36 -12 38
rect 36 44 38 46
rect 50 44 52 46
rect 26 36 28 38
rect 141 44 143 46
rect 155 44 157 46
rect 66 31 68 33
rect 131 36 133 38
rect 171 31 173 33
<< ndifct0 >>
rect -11 27 -9 29
rect -20 14 -18 16
rect 50 27 52 29
rect 39 20 41 22
rect 64 19 66 21
rect -1 14 1 16
rect 76 22 78 24
rect 155 27 157 29
rect 144 20 146 22
rect 169 19 171 21
rect 181 22 183 24
<< ndifct1 >>
rect -31 27 -29 29
rect 9 22 11 24
rect 86 20 88 22
rect 20 10 22 12
rect 114 22 116 24
rect 104 10 106 12
rect 191 20 193 22
rect 125 10 127 12
rect 209 10 211 12
<< ntiect1 >>
rect -30 70 -28 72
rect 10 70 12 72
rect 84 70 86 72
rect 115 70 117 72
rect 189 70 191 72
<< ptiect1 >>
rect -30 10 -28 12
rect 10 10 12 12
rect 51 10 53 12
rect 115 10 117 12
rect 156 10 158 12
<< pdifct0 >>
rect -20 67 -18 69
rect -1 60 1 62
rect 19 58 21 60
rect 29 60 31 62
rect 29 53 31 55
rect 39 60 41 62
rect 58 46 60 48
rect 68 67 70 69
rect 68 60 70 62
rect 84 53 86 55
rect 84 46 86 48
rect 104 61 106 63
rect 124 58 126 60
rect 134 60 136 62
rect 134 53 136 55
rect 144 60 146 62
rect 163 46 165 48
rect 173 67 175 69
rect 173 60 175 62
rect 189 53 191 55
rect 189 46 191 48
rect 209 61 211 63
<< pdifct1 >>
rect -31 57 -29 59
rect -31 50 -29 52
rect 9 53 11 55
rect 9 46 11 48
rect 94 53 96 55
rect 114 53 116 55
rect 114 46 116 48
rect 199 53 201 55
<< alu0 >>
rect -22 67 -20 69
rect -18 67 -16 69
rect -22 66 -16 67
rect -14 62 3 63
rect -14 60 -1 62
rect 1 60 3 62
rect -14 59 3 60
rect 17 60 23 69
rect -29 48 -28 59
rect -14 55 -10 59
rect 17 58 19 60
rect 21 58 23 60
rect 17 57 23 58
rect 28 62 32 64
rect 28 60 29 62
rect 31 60 32 62
rect -25 51 -10 55
rect -25 38 -21 51
rect 28 55 32 60
rect 37 62 43 69
rect 67 67 68 69
rect 70 67 71 69
rect 37 60 39 62
rect 41 60 43 62
rect 37 59 43 60
rect 67 62 71 67
rect 67 60 68 62
rect 70 60 71 62
rect 67 58 71 60
rect 75 63 108 64
rect 75 61 104 63
rect 106 61 108 63
rect 75 60 108 61
rect 122 60 128 69
rect 28 54 29 55
rect 15 53 29 54
rect 31 53 32 55
rect 15 50 32 53
rect -6 42 0 43
rect -25 36 -24 38
rect -22 36 -21 38
rect -25 30 -21 36
rect -25 29 -7 30
rect -25 27 -11 29
rect -9 27 -7 29
rect -25 26 -7 27
rect 15 38 19 50
rect 75 49 79 60
rect 122 58 124 60
rect 126 58 128 60
rect 122 57 128 58
rect 133 62 137 64
rect 133 60 134 62
rect 136 60 137 62
rect 56 48 79 49
rect 56 46 58 48
rect 60 46 79 48
rect 56 45 79 46
rect 56 39 60 45
rect 15 36 16 38
rect 18 36 19 38
rect 15 31 19 36
rect 15 27 27 31
rect 11 24 12 26
rect 23 23 27 27
rect 49 35 60 39
rect 49 29 53 35
rect 75 39 79 45
rect 83 55 87 57
rect 83 53 84 55
rect 86 53 87 55
rect 83 48 87 53
rect 83 46 84 48
rect 86 47 87 48
rect 86 46 99 47
rect 83 43 99 46
rect 95 41 99 43
rect 95 39 100 41
rect 75 38 91 39
rect 75 36 87 38
rect 89 36 91 38
rect 75 35 91 36
rect 95 37 97 39
rect 99 37 100 39
rect 95 35 100 37
rect 49 27 50 29
rect 52 27 53 29
rect 49 25 53 27
rect 95 31 99 35
rect 75 27 99 31
rect 75 24 79 27
rect 23 22 43 23
rect 75 22 76 24
rect 78 22 79 24
rect 23 20 39 22
rect 41 20 43 22
rect 23 19 43 20
rect 62 21 68 22
rect 62 19 64 21
rect 66 19 68 21
rect 75 20 79 22
rect 133 55 137 60
rect 142 62 148 69
rect 172 67 173 69
rect 175 67 176 69
rect 142 60 144 62
rect 146 60 148 62
rect 142 59 148 60
rect 172 62 176 67
rect 172 60 173 62
rect 175 60 176 62
rect 172 58 176 60
rect 180 63 213 64
rect 180 61 209 63
rect 211 61 213 63
rect 180 60 213 61
rect 133 54 134 55
rect 120 53 134 54
rect 136 53 137 55
rect 120 50 137 53
rect 120 38 124 50
rect 180 49 184 60
rect 161 48 184 49
rect 161 46 163 48
rect 165 46 184 48
rect 161 45 184 46
rect 161 39 165 45
rect 120 36 121 38
rect 123 36 124 38
rect 120 31 124 36
rect 120 27 132 31
rect 116 24 117 26
rect -22 16 -16 17
rect -22 14 -20 16
rect -18 14 -16 16
rect -22 13 -16 14
rect -3 16 3 17
rect -3 14 -1 16
rect 1 14 3 16
rect -3 13 3 14
rect 62 13 68 19
rect 128 23 132 27
rect 154 35 165 39
rect 154 29 158 35
rect 180 39 184 45
rect 188 55 192 57
rect 188 53 189 55
rect 191 53 192 55
rect 188 48 192 53
rect 188 46 189 48
rect 191 47 192 48
rect 191 46 204 47
rect 188 43 204 46
rect 200 41 204 43
rect 200 39 205 41
rect 180 38 196 39
rect 180 36 192 38
rect 194 36 196 38
rect 180 35 196 36
rect 200 37 202 39
rect 204 37 205 39
rect 200 35 205 37
rect 154 27 155 29
rect 157 27 158 29
rect 154 25 158 27
rect 200 31 204 35
rect 180 27 204 31
rect 180 24 184 27
rect 128 22 148 23
rect 180 22 181 24
rect 183 22 184 24
rect 128 20 144 22
rect 146 20 148 22
rect 128 19 148 20
rect 167 21 173 22
rect 167 19 169 21
rect 171 19 173 21
rect 180 20 184 22
rect 167 13 173 19
<< via1 >>
rect 0 53 2 55
rect 32 27 34 29
rect 59 27 61 29
rect 105 27 107 29
rect 114 53 116 55
rect 137 27 139 29
rect 164 27 166 29
<< labels >>
rlabel alu1 58 61 58 61 6 b
rlabel alu1 49 73 49 73 1 Vdd
rlabel alu1 33 33 33 33 6 a
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 41 53 41 53 6 b
rlabel alu1 47 8 47 8 1 Vss
rlabel alu1 67 36 67 36 1 a
rlabel alu1 154 73 154 73 1 Vdd
rlabel alu1 211 40 211 40 1 sum
rlabel alu1 130 73 130 73 6 vdd
rlabel alu1 152 8 152 8 1 Vss
rlabel alu1 146 53 146 53 1 cin
rlabel alu1 139 34 139 34 1 s0
rlabel alu1 106 40 106 40 1 s0
rlabel alu1 171 28 171 28 1 s0
rlabel alu1 114 34 114 34 1 c0
rlabel alu1 9 35 9 35 1 c1
rlabel alu1 -15 73 -15 73 6 vdd
rlabel alu1 1 29 1 29 1 c1
rlabel alu1 1 53 1 53 1 c0
rlabel alu1 -31 44 -31 44 1 cout
<< end >>
