magic
tech scmos
timestamp 1607610918
<< ab >>
rect 4 136 68 154
rect 74 146 142 154
rect -1 131 68 136
rect 78 131 142 146
rect 6 109 68 131
rect 6 108 11 109
rect 13 108 68 109
rect 6 90 68 108
rect 80 124 142 131
rect 80 119 147 124
rect 80 90 142 119
rect 4 82 68 90
rect 78 82 142 90
rect 144 82 147 90
rect 2 77 70 82
rect 2 69 22 77
rect 3 5 22 13
rect 24 5 64 77
rect 66 69 70 77
rect 76 77 147 82
rect 76 69 96 77
rect 66 5 96 13
rect 98 5 138 77
rect 140 69 147 77
rect 102 -33 142 -4
rect 102 -38 147 -33
rect 102 -45 142 -38
rect 104 -49 142 -45
rect 97 -76 101 -68
rect 102 -76 142 -49
<< nwell >>
rect -1 114 147 159
rect -1 5 147 45
rect 63 -44 147 5
<< pwell >>
rect -1 45 147 114
rect 63 -81 147 -44
<< poly >>
rect 21 148 23 152
rect 6 123 12 125
rect 6 121 8 123
rect 10 121 12 123
rect 57 148 59 152
rect 95 148 97 152
rect 37 139 39 143
rect 47 139 49 143
rect 80 123 86 125
rect 80 121 82 123
rect 84 121 86 123
rect 131 148 133 152
rect 111 139 113 143
rect 121 139 123 143
rect 6 119 12 121
rect 10 118 12 119
rect 21 118 23 121
rect 37 118 39 121
rect 10 116 23 118
rect 29 116 39 118
rect 47 117 49 121
rect 57 118 59 121
rect 80 119 86 121
rect 13 108 15 116
rect 29 112 31 116
rect 22 110 31 112
rect 43 115 49 117
rect 43 113 45 115
rect 47 113 49 115
rect 43 111 49 113
rect 53 116 59 118
rect 84 118 86 119
rect 95 118 97 121
rect 111 118 113 121
rect 84 116 97 118
rect 103 116 113 118
rect 121 117 123 121
rect 131 118 133 121
rect 53 114 55 116
rect 57 114 59 116
rect 53 112 59 114
rect 22 108 24 110
rect 26 108 31 110
rect 22 106 31 108
rect 47 108 49 111
rect 29 103 31 106
rect 39 103 41 107
rect 47 106 51 108
rect 49 103 51 106
rect 56 103 58 112
rect 87 108 89 116
rect 103 112 105 116
rect 96 110 105 112
rect 117 115 123 117
rect 117 113 119 115
rect 121 113 123 115
rect 117 111 123 113
rect 127 116 133 118
rect 127 114 129 116
rect 131 114 133 116
rect 127 112 133 114
rect 96 108 98 110
rect 100 108 105 110
rect 13 96 15 99
rect 13 94 18 96
rect 16 86 18 94
rect 29 90 31 94
rect 39 86 41 94
rect 96 106 105 108
rect 121 108 123 111
rect 103 103 105 106
rect 113 103 115 107
rect 121 106 125 108
rect 123 103 125 106
rect 130 103 132 112
rect 87 96 89 99
rect 87 94 92 96
rect 49 86 51 91
rect 56 86 58 91
rect 16 84 41 86
rect 90 86 92 94
rect 103 90 105 94
rect 113 86 115 94
rect 123 86 125 91
rect 130 86 132 91
rect 90 84 115 86
rect 33 64 35 69
rect 40 64 42 69
rect 53 62 55 66
rect 107 64 109 69
rect 114 64 116 69
rect 127 62 129 66
rect 33 40 35 53
rect 40 48 42 53
rect 53 48 55 53
rect 39 46 45 48
rect 39 44 41 46
rect 43 44 45 46
rect 39 42 45 44
rect 49 46 55 48
rect 49 44 51 46
rect 53 44 55 46
rect 49 42 55 44
rect 29 38 35 40
rect 29 36 31 38
rect 33 36 35 38
rect 29 34 35 36
rect 33 31 35 34
rect 43 31 45 42
rect 53 38 55 42
rect 107 40 109 53
rect 114 48 116 53
rect 127 48 129 53
rect 113 46 119 48
rect 113 44 115 46
rect 117 44 119 46
rect 113 42 119 44
rect 123 46 129 48
rect 123 44 125 46
rect 127 44 129 46
rect 123 42 129 44
rect 103 38 109 40
rect 103 36 105 38
rect 107 36 109 38
rect 103 34 109 36
rect 107 31 109 34
rect 117 31 119 42
rect 127 38 129 42
rect 33 13 35 18
rect 43 13 45 18
rect 53 16 55 20
rect 107 13 109 18
rect 117 13 119 18
rect 127 16 129 20
rect 111 -10 113 -6
rect 118 -10 120 -6
rect 131 -20 133 -15
rect 111 -34 113 -31
rect 107 -36 113 -34
rect 107 -38 109 -36
rect 111 -38 113 -36
rect 107 -40 113 -38
rect 111 -50 113 -40
rect 118 -41 120 -31
rect 131 -41 133 -38
rect 117 -43 123 -41
rect 117 -45 119 -43
rect 121 -45 123 -43
rect 117 -47 123 -45
rect 127 -43 133 -41
rect 127 -45 129 -43
rect 131 -45 133 -43
rect 127 -47 133 -45
rect 121 -50 123 -47
rect 131 -50 133 -47
rect 111 -61 113 -56
rect 121 -61 123 -56
rect 131 -64 133 -59
<< ndif >>
rect 6 102 13 108
rect 8 99 13 102
rect 15 103 20 108
rect 80 106 87 108
rect 80 104 82 106
rect 84 104 87 106
rect 15 99 29 103
rect 20 98 29 99
rect 20 96 22 98
rect 24 96 29 98
rect 20 94 29 96
rect 31 101 39 103
rect 31 99 34 101
rect 36 99 39 101
rect 31 94 39 99
rect 41 99 49 103
rect 41 97 44 99
rect 46 97 49 99
rect 41 94 49 97
rect 44 91 49 94
rect 51 91 56 103
rect 58 91 66 103
rect 80 102 87 104
rect 82 99 87 102
rect 89 103 94 108
rect 89 99 103 103
rect 94 98 103 99
rect 94 96 96 98
rect 98 96 103 98
rect 94 94 103 96
rect 105 101 113 103
rect 105 99 108 101
rect 110 99 113 101
rect 105 94 113 99
rect 115 99 123 103
rect 115 97 118 99
rect 120 97 123 99
rect 115 94 123 97
rect 60 89 66 91
rect 60 87 62 89
rect 64 87 66 89
rect 60 85 66 87
rect 118 91 123 94
rect 125 91 130 103
rect 132 91 140 103
rect 134 89 140 91
rect 134 87 136 89
rect 138 87 140 89
rect 134 85 140 87
rect 44 72 51 74
rect 44 70 47 72
rect 49 70 51 72
rect 44 64 51 70
rect 118 72 125 74
rect 118 70 121 72
rect 123 70 125 72
rect 26 62 33 64
rect 26 60 28 62
rect 30 60 33 62
rect 26 58 33 60
rect 28 53 33 58
rect 35 53 40 64
rect 42 62 51 64
rect 118 64 125 70
rect 100 62 107 64
rect 42 53 53 62
rect 55 60 62 62
rect 55 58 58 60
rect 60 58 62 60
rect 100 60 102 62
rect 104 60 107 62
rect 100 58 107 60
rect 55 56 62 58
rect 55 53 60 56
rect 102 53 107 58
rect 109 53 114 64
rect 116 62 125 64
rect 116 53 127 62
rect 129 60 136 62
rect 129 58 132 60
rect 134 58 136 60
rect 129 56 136 58
rect 129 53 134 56
rect 104 -56 111 -50
rect 113 -52 121 -50
rect 113 -54 116 -52
rect 118 -54 121 -52
rect 113 -56 121 -54
rect 123 -56 131 -50
rect 104 -63 109 -56
rect 125 -59 131 -56
rect 133 -52 140 -50
rect 133 -54 136 -52
rect 138 -54 140 -52
rect 133 -56 140 -54
rect 133 -59 138 -56
rect 125 -63 129 -59
rect 104 -65 110 -63
rect 104 -67 106 -65
rect 108 -67 110 -65
rect 104 -69 110 -67
rect 123 -65 129 -63
rect 123 -67 125 -65
rect 127 -67 129 -65
rect 123 -69 129 -67
<< pdif >>
rect 16 127 21 148
rect 14 125 21 127
rect 14 123 16 125
rect 18 123 21 125
rect 14 121 21 123
rect 23 146 35 148
rect 23 144 26 146
rect 28 144 35 146
rect 23 139 35 144
rect 52 139 57 148
rect 23 137 26 139
rect 28 137 37 139
rect 23 121 37 137
rect 39 132 47 139
rect 39 130 42 132
rect 44 130 47 132
rect 39 125 47 130
rect 39 123 42 125
rect 44 123 47 125
rect 39 121 47 123
rect 49 132 57 139
rect 49 130 52 132
rect 54 130 57 132
rect 49 121 57 130
rect 59 142 64 148
rect 59 140 66 142
rect 59 138 62 140
rect 64 138 66 140
rect 59 136 66 138
rect 59 121 64 136
rect 90 127 95 148
rect 88 125 95 127
rect 88 123 90 125
rect 92 123 95 125
rect 88 121 95 123
rect 97 146 109 148
rect 97 144 100 146
rect 102 144 109 146
rect 97 139 109 144
rect 126 139 131 148
rect 97 137 100 139
rect 102 137 111 139
rect 97 121 111 137
rect 113 132 121 139
rect 113 130 116 132
rect 118 130 121 132
rect 113 125 121 130
rect 113 123 116 125
rect 118 123 121 125
rect 113 121 121 123
rect 123 132 131 139
rect 123 130 126 132
rect 128 130 131 132
rect 123 121 131 130
rect 133 142 138 148
rect 133 140 140 142
rect 133 138 136 140
rect 138 138 140 140
rect 133 136 140 138
rect 133 121 138 136
rect 47 31 53 38
rect 26 22 33 31
rect 26 20 28 22
rect 30 20 33 22
rect 26 18 33 20
rect 35 29 43 31
rect 35 27 38 29
rect 40 27 43 29
rect 35 22 43 27
rect 35 20 38 22
rect 40 20 43 22
rect 35 18 43 20
rect 45 24 53 31
rect 45 22 48 24
rect 50 22 53 24
rect 45 20 53 22
rect 55 36 62 38
rect 55 34 58 36
rect 60 34 62 36
rect 55 29 62 34
rect 121 31 127 38
rect 55 27 58 29
rect 60 27 62 29
rect 55 25 62 27
rect 55 20 60 25
rect 100 22 107 31
rect 100 20 102 22
rect 104 20 107 22
rect 45 18 51 20
rect 100 18 107 20
rect 109 29 117 31
rect 109 27 112 29
rect 114 27 117 29
rect 109 22 117 27
rect 109 20 112 22
rect 114 20 117 22
rect 109 18 117 20
rect 119 24 127 31
rect 119 22 122 24
rect 124 22 127 24
rect 119 20 127 22
rect 129 36 136 38
rect 129 34 132 36
rect 134 34 136 36
rect 129 29 136 34
rect 129 27 132 29
rect 134 27 136 29
rect 129 25 136 27
rect 129 20 134 25
rect 119 18 125 20
rect 106 -17 111 -10
rect 104 -19 111 -17
rect 104 -21 106 -19
rect 108 -21 111 -19
rect 104 -23 111 -21
rect 106 -31 111 -23
rect 113 -31 118 -10
rect 120 -12 129 -10
rect 120 -14 125 -12
rect 127 -14 129 -12
rect 120 -20 129 -14
rect 120 -31 131 -20
rect 123 -38 131 -31
rect 133 -22 140 -20
rect 133 -24 136 -22
rect 138 -24 140 -22
rect 133 -29 140 -24
rect 133 -31 136 -29
rect 138 -31 140 -29
rect 133 -33 140 -31
rect 133 -38 138 -33
<< alu1 >>
rect 2 149 144 154
rect 2 147 42 149
rect 44 147 116 149
rect 118 147 144 149
rect 2 146 144 147
rect 6 136 18 141
rect -1 135 18 136
rect -1 131 11 135
rect 6 129 11 131
rect 6 127 7 129
rect 9 127 11 129
rect 6 123 11 127
rect 80 135 92 141
rect 6 121 8 123
rect 10 121 11 123
rect 6 119 11 121
rect 22 110 27 117
rect 80 133 85 135
rect 50 132 85 133
rect 50 130 52 132
rect 54 130 85 132
rect 50 129 85 130
rect 50 128 81 129
rect 62 127 81 128
rect 83 127 85 129
rect 22 109 24 110
rect 14 108 24 109
rect 26 108 27 110
rect 14 106 27 108
rect 14 104 18 106
rect 20 104 27 106
rect 14 103 27 104
rect 62 100 66 127
rect 80 123 85 127
rect 80 121 82 123
rect 84 121 85 123
rect 80 119 85 121
rect 96 110 101 117
rect 124 132 140 133
rect 124 130 126 132
rect 128 130 140 132
rect 124 128 140 130
rect 136 124 140 128
rect 136 119 147 124
rect 96 109 98 110
rect 88 108 98 109
rect 100 108 101 110
rect 88 106 101 108
rect 88 104 92 106
rect 94 104 101 106
rect 88 103 101 104
rect 42 99 66 100
rect 136 100 140 119
rect 42 97 44 99
rect 46 97 66 99
rect 42 96 66 97
rect 116 99 140 100
rect 116 97 118 99
rect 120 97 140 99
rect 116 96 140 97
rect 2 89 147 90
rect 2 87 9 89
rect 11 87 62 89
rect 64 87 83 89
rect 85 87 136 89
rect 138 87 147 89
rect 2 72 147 87
rect 2 70 47 72
rect 49 70 57 72
rect 59 70 121 72
rect 123 70 131 72
rect 133 70 147 72
rect 2 69 147 70
rect 33 48 38 56
rect 50 60 62 64
rect 50 58 58 60
rect 60 58 62 60
rect 33 46 34 48
rect 36 47 38 48
rect 36 46 47 47
rect 33 44 41 46
rect 43 44 47 46
rect 33 43 47 44
rect 26 38 39 39
rect 26 36 31 38
rect 33 36 39 38
rect 26 35 39 36
rect 26 34 30 35
rect 26 32 27 34
rect 29 32 30 34
rect 58 48 62 58
rect 58 46 59 48
rect 61 46 62 48
rect 58 38 62 46
rect 107 48 112 56
rect 124 60 136 64
rect 124 58 132 60
rect 134 58 136 60
rect 107 46 108 48
rect 110 47 112 48
rect 110 46 121 47
rect 107 44 115 46
rect 117 44 121 46
rect 107 43 121 44
rect 26 26 30 32
rect 57 36 62 38
rect 57 34 58 36
rect 60 34 62 36
rect 57 29 62 34
rect 57 27 58 29
rect 60 27 62 29
rect 57 21 62 27
rect 100 38 113 39
rect 100 36 105 38
rect 107 36 113 38
rect 100 35 113 36
rect 100 34 104 35
rect 100 32 101 34
rect 103 32 104 34
rect 132 49 136 58
rect 132 47 133 49
rect 135 47 136 49
rect 132 38 136 47
rect 100 26 104 32
rect 131 36 136 38
rect 131 34 132 36
rect 134 34 136 36
rect 131 29 136 34
rect 131 27 132 29
rect 134 27 136 29
rect 131 25 136 27
rect 3 12 147 13
rect 3 10 57 12
rect 59 10 131 12
rect 133 10 147 12
rect 3 5 147 10
rect 63 -9 144 -4
rect 63 -11 135 -9
rect 137 -11 144 -9
rect 63 -12 144 -11
rect 136 -18 140 -17
rect 127 -22 140 -18
rect 104 -34 108 -25
rect 104 -35 125 -34
rect 104 -37 105 -35
rect 107 -36 125 -35
rect 107 -37 109 -36
rect 104 -38 109 -37
rect 111 -38 125 -36
rect 104 -43 125 -42
rect 104 -45 105 -43
rect 107 -45 119 -43
rect 121 -45 125 -43
rect 104 -46 125 -45
rect 138 -24 140 -22
rect 136 -29 140 -24
rect 138 -31 140 -29
rect 136 -33 140 -31
rect 104 -55 108 -46
rect 136 -38 147 -33
rect 136 -50 140 -38
rect 135 -52 140 -50
rect 135 -54 136 -52
rect 138 -54 140 -52
rect 135 -56 140 -54
rect 97 -69 144 -68
rect 97 -71 135 -69
rect 137 -71 144 -69
rect 97 -76 144 -71
<< alu2 >>
rect 6 129 11 131
rect 6 127 7 129
rect 9 127 11 129
rect 6 35 11 127
rect 80 129 85 131
rect 80 127 81 129
rect 83 127 85 129
rect 17 106 21 109
rect 17 104 18 106
rect 20 104 21 106
rect 17 50 21 104
rect 17 48 38 50
rect 17 46 34 48
rect 36 46 38 48
rect 17 45 38 46
rect 58 48 72 49
rect 58 46 59 48
rect 61 46 72 48
rect 58 45 72 46
rect 6 34 30 35
rect 6 32 27 34
rect 29 32 30 34
rect 6 31 30 32
rect 67 -34 72 45
rect 80 35 85 127
rect 91 106 95 109
rect 91 104 92 106
rect 94 104 95 106
rect 91 50 95 104
rect 91 48 112 50
rect 91 46 108 48
rect 110 46 112 48
rect 132 49 144 50
rect 132 47 133 49
rect 135 47 144 49
rect 132 46 144 47
rect 91 45 112 46
rect 80 34 104 35
rect 80 32 101 34
rect 103 32 104 34
rect 80 31 104 32
rect 67 -35 108 -34
rect 67 -37 105 -35
rect 107 -37 108 -35
rect 67 -38 108 -37
rect 96 -43 108 -42
rect 96 -45 105 -43
rect 107 -45 108 -43
rect 96 -46 108 -45
rect 96 -61 100 -46
rect 139 -61 144 46
rect 96 -66 144 -61
<< ptie >>
rect 7 89 13 91
rect 7 87 9 89
rect 11 87 13 89
rect 7 85 13 87
rect 81 89 87 91
rect 81 87 83 89
rect 85 87 87 89
rect 81 85 87 87
rect 55 72 61 74
rect 55 70 57 72
rect 59 70 61 72
rect 55 68 61 70
rect 129 72 135 74
rect 129 70 131 72
rect 133 70 135 72
rect 129 68 135 70
rect 133 -69 139 -67
rect 133 -71 135 -69
rect 137 -71 139 -69
rect 133 -73 139 -71
<< ntie >>
rect 40 149 46 151
rect 40 147 42 149
rect 44 147 46 149
rect 114 149 120 151
rect 40 145 46 147
rect 114 147 116 149
rect 118 147 120 149
rect 114 145 120 147
rect 55 12 61 14
rect 55 10 57 12
rect 59 10 61 12
rect 55 8 61 10
rect 129 12 135 14
rect 129 10 131 12
rect 133 10 135 12
rect 129 8 135 10
rect 133 -9 139 -7
rect 133 -11 135 -9
rect 137 -11 139 -9
rect 133 -13 139 -11
<< nmos >>
rect 13 99 15 108
rect 29 94 31 103
rect 39 94 41 103
rect 49 91 51 103
rect 56 91 58 103
rect 87 99 89 108
rect 103 94 105 103
rect 113 94 115 103
rect 123 91 125 103
rect 130 91 132 103
rect 33 53 35 64
rect 40 53 42 64
rect 53 53 55 62
rect 107 53 109 64
rect 114 53 116 64
rect 127 53 129 62
rect 111 -56 113 -50
rect 121 -56 123 -50
rect 131 -59 133 -50
<< pmos >>
rect 21 121 23 148
rect 37 121 39 139
rect 47 121 49 139
rect 57 121 59 148
rect 95 121 97 148
rect 111 121 113 139
rect 121 121 123 139
rect 131 121 133 148
rect 33 18 35 31
rect 43 18 45 31
rect 53 20 55 38
rect 107 18 109 31
rect 117 18 119 31
rect 127 20 129 38
rect 111 -31 113 -10
rect 118 -31 120 -10
rect 131 -38 133 -20
<< polyct0 >>
rect 45 113 47 115
rect 55 114 57 116
rect 119 113 121 115
rect 129 114 131 116
rect 51 44 53 46
rect 125 44 127 46
rect 129 -45 131 -43
<< polyct1 >>
rect 8 121 10 123
rect 82 121 84 123
rect 24 108 26 110
rect 98 108 100 110
rect 41 44 43 46
rect 31 36 33 38
rect 115 44 117 46
rect 105 36 107 38
rect 109 -38 111 -36
rect 119 -45 121 -43
<< ndifct0 >>
rect 82 104 84 106
rect 22 96 24 98
rect 34 99 36 101
rect 96 96 98 98
rect 108 99 110 101
rect 28 60 30 62
rect 102 60 104 62
rect 116 -54 118 -52
rect 106 -67 108 -65
rect 125 -67 127 -65
<< ndifct1 >>
rect 44 97 46 99
rect 118 97 120 99
rect 62 87 64 89
rect 136 87 138 89
rect 47 70 49 72
rect 121 70 123 72
rect 58 58 60 60
rect 132 58 134 60
rect 136 -54 138 -52
<< ntiect1 >>
rect 42 147 44 149
rect 116 147 118 149
rect 57 10 59 12
rect 131 10 133 12
rect 135 -11 137 -9
<< ptiect1 >>
rect 9 87 11 89
rect 83 87 85 89
rect 57 70 59 72
rect 131 70 133 72
rect 135 -71 137 -69
<< pdifct0 >>
rect 16 123 18 125
rect 26 144 28 146
rect 26 137 28 139
rect 42 130 44 132
rect 42 123 44 125
rect 62 138 64 140
rect 90 123 92 125
rect 100 144 102 146
rect 100 137 102 139
rect 116 130 118 132
rect 116 123 118 125
rect 136 138 138 140
rect 28 20 30 22
rect 38 27 40 29
rect 38 20 40 22
rect 48 22 50 24
rect 102 20 104 22
rect 112 27 114 29
rect 112 20 114 22
rect 122 22 124 24
rect 106 -21 108 -19
rect 125 -14 127 -12
<< pdifct1 >>
rect 52 130 54 132
rect 126 130 128 132
rect 58 34 60 36
rect 58 27 60 29
rect 132 34 134 36
rect 132 27 134 29
rect 136 -24 138 -22
rect 136 -31 138 -29
<< alu0 >>
rect 25 144 26 146
rect 28 144 29 146
rect 25 139 29 144
rect 99 144 100 146
rect 102 144 103 146
rect 25 137 26 139
rect 28 137 29 139
rect 25 135 29 137
rect 33 140 66 141
rect 33 138 62 140
rect 64 138 66 140
rect 33 137 66 138
rect 33 126 37 137
rect 99 139 103 144
rect 99 137 100 139
rect 102 137 103 139
rect 99 135 103 137
rect 107 140 140 141
rect 107 138 136 140
rect 138 138 140 140
rect 107 137 140 138
rect 14 125 37 126
rect 14 123 16 125
rect 18 123 37 125
rect 14 122 37 123
rect 14 116 18 122
rect 7 112 18 116
rect 7 102 11 112
rect 33 116 37 122
rect 41 132 45 134
rect 41 130 42 132
rect 44 130 45 132
rect 41 125 45 130
rect 41 123 42 125
rect 44 124 45 125
rect 44 123 57 124
rect 41 120 57 123
rect 53 118 57 120
rect 53 116 58 118
rect 33 115 49 116
rect 33 113 45 115
rect 47 113 49 115
rect 33 112 49 113
rect 53 114 55 116
rect 57 114 58 116
rect 53 112 58 114
rect 53 108 57 112
rect 33 104 57 108
rect 33 101 37 104
rect 33 99 34 101
rect 36 99 37 101
rect 107 126 111 137
rect 88 125 111 126
rect 88 123 90 125
rect 92 123 111 125
rect 88 122 111 123
rect 88 116 92 122
rect 81 112 92 116
rect 81 106 85 112
rect 107 116 111 122
rect 115 132 119 134
rect 115 130 116 132
rect 118 130 119 132
rect 115 125 119 130
rect 115 123 116 125
rect 118 124 119 125
rect 118 123 131 124
rect 115 120 131 123
rect 127 118 131 120
rect 127 116 132 118
rect 107 115 123 116
rect 107 113 119 115
rect 121 113 123 115
rect 107 112 123 113
rect 127 114 129 116
rect 131 114 132 116
rect 127 112 132 114
rect 81 104 82 106
rect 84 104 85 106
rect 81 102 85 104
rect 127 108 131 112
rect 107 104 131 108
rect 20 98 26 99
rect 20 96 22 98
rect 24 96 26 98
rect 33 97 37 99
rect 107 101 111 104
rect 107 99 108 101
rect 110 99 111 101
rect 94 98 100 99
rect 94 96 96 98
rect 98 96 100 98
rect 107 97 111 99
rect 20 90 26 96
rect 94 90 100 96
rect 26 62 46 63
rect 26 60 28 62
rect 30 60 46 62
rect 26 59 46 60
rect 42 55 46 59
rect 100 62 120 63
rect 100 60 102 62
rect 104 60 120 62
rect 100 59 120 60
rect 57 56 58 58
rect 42 51 54 55
rect 50 46 54 51
rect 50 44 51 46
rect 53 44 54 46
rect 50 32 54 44
rect 116 55 120 59
rect 131 56 132 58
rect 116 51 128 55
rect 124 46 128 51
rect 124 44 125 46
rect 127 44 128 46
rect 37 29 54 32
rect 37 27 38 29
rect 40 28 54 29
rect 40 27 41 28
rect 26 22 32 23
rect 26 20 28 22
rect 30 20 32 22
rect 26 13 32 20
rect 37 22 41 27
rect 37 20 38 22
rect 40 20 41 22
rect 37 18 41 20
rect 46 24 52 25
rect 46 22 48 24
rect 50 22 52 24
rect 46 13 52 22
rect 124 32 128 44
rect 111 29 128 32
rect 111 27 112 29
rect 114 28 128 29
rect 114 27 115 28
rect 100 22 106 23
rect 100 20 102 22
rect 104 20 106 22
rect 100 13 106 20
rect 111 22 115 27
rect 111 20 112 22
rect 114 20 115 22
rect 111 18 115 20
rect 120 24 126 25
rect 120 22 122 24
rect 124 22 126 24
rect 120 13 126 22
rect 123 -14 125 -12
rect 127 -14 129 -12
rect 123 -15 129 -14
rect 104 -19 121 -18
rect 104 -21 106 -19
rect 108 -21 121 -19
rect 104 -22 121 -21
rect 117 -26 121 -22
rect 117 -30 132 -26
rect 107 -39 113 -38
rect 128 -43 132 -30
rect 135 -33 136 -22
rect 128 -45 129 -43
rect 131 -45 132 -43
rect 128 -51 132 -45
rect 114 -52 132 -51
rect 114 -54 116 -52
rect 118 -54 132 -52
rect 114 -55 132 -54
rect 104 -65 110 -64
rect 104 -67 106 -65
rect 108 -67 110 -65
rect 104 -68 110 -67
rect 123 -65 129 -64
rect 123 -67 125 -65
rect 127 -67 129 -65
rect 123 -68 129 -67
<< via1 >>
rect 7 127 9 129
rect 81 127 83 129
rect 18 104 20 106
rect 92 104 94 106
rect 34 46 36 48
rect 27 32 29 34
rect 59 46 61 48
rect 108 46 110 48
rect 101 32 103 34
rect 133 47 135 49
rect 105 -37 107 -35
rect 105 -45 107 -43
<< labels >>
rlabel alu1 8 130 8 130 6 b
rlabel alu1 36 150 36 150 6 vdd
rlabel alu1 28 29 28 29 2 b
rlabel alu1 44 9 44 9 2 vdd
rlabel alu1 36 49 36 49 2 a
rlabel alu1 138 119 138 119 1 sum
rlabel alu1 64 119 64 120 1 s1
rlabel alu1 82 131 82 132 1 s1
rlabel alu1 122 -72 122 -72 4 vss
rlabel alu1 122 -8 122 -8 4 vdd
rlabel alu1 138 -36 138 -36 5 cout
rlabel alu2 136 46 136 50 1 cout2
rlabel alu2 62 45 62 49 1 cout1
rlabel alu1 140 119 140 123 1 sum
rlabel alu1 140 -38 140 -34 1 cout
rlabel alu1 72 78 72 79 1 vss
rlabel alu1 0 131 0 136 3 b
rlabel alu1 23 109 23 109 1 a
rlabel via1 93 105 93 105 1 cin
rlabel via1 105 -45 105 -45 1 cout2
rlabel via1 109 47 109 47 1 cin
<< end >>
