magic
tech scmos
timestamp 1607768000
<< ab >>
rect 5 5 45 77
rect 47 69 52 77
rect 54 69 158 77
rect 54 37 94 69
rect 95 37 158 69
rect 54 5 158 37
rect 168 69 272 77
rect 273 69 275 77
rect 168 37 208 69
rect 209 37 272 69
rect 168 5 272 37
rect 273 5 277 13
rect 279 5 319 77
rect 320 69 384 77
rect 323 13 384 69
rect 320 5 384 13
rect 388 5 452 77
rect 456 5 519 77
rect 521 69 561 77
rect 562 69 627 77
rect 628 69 633 77
rect 522 13 561 69
rect 564 13 627 69
rect 521 5 561 13
rect 563 5 633 13
rect 89 0 95 5
rect 203 0 209 5
<< nwell >>
rect 0 37 633 82
<< pwell >>
rect 0 0 633 37
<< poly >>
rect 27 71 29 75
rect 34 71 36 75
rect 14 61 16 66
rect 111 71 113 75
rect 63 62 65 66
rect 73 64 75 69
rect 83 64 85 69
rect 14 40 16 43
rect 27 40 29 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 31 16 34
rect 24 31 26 34
rect 34 31 36 41
rect 63 40 65 44
rect 73 40 75 51
rect 83 48 85 51
rect 83 46 89 48
rect 83 44 85 46
rect 87 44 89 46
rect 83 42 89 44
rect 96 46 102 48
rect 96 44 98 46
rect 100 44 102 46
rect 147 71 149 75
rect 127 62 129 66
rect 137 62 139 66
rect 225 71 227 75
rect 177 62 179 66
rect 187 64 189 69
rect 197 64 199 69
rect 96 42 102 44
rect 63 38 69 40
rect 63 36 65 38
rect 67 36 69 38
rect 63 34 69 36
rect 73 38 79 40
rect 73 36 75 38
rect 77 36 79 38
rect 73 34 79 36
rect 63 29 65 34
rect 76 29 78 34
rect 83 29 85 42
rect 100 41 102 42
rect 111 41 113 44
rect 127 41 129 44
rect 100 39 113 41
rect 119 39 129 41
rect 137 40 139 44
rect 147 41 149 44
rect 103 31 105 39
rect 119 35 121 39
rect 112 33 121 35
rect 133 38 139 40
rect 133 36 135 38
rect 137 36 139 38
rect 133 34 139 36
rect 143 39 149 41
rect 143 37 145 39
rect 147 37 149 39
rect 143 35 149 37
rect 177 40 179 44
rect 187 40 189 51
rect 197 48 199 51
rect 197 46 203 48
rect 197 44 199 46
rect 201 44 203 46
rect 197 42 203 44
rect 210 46 216 48
rect 210 44 212 46
rect 214 44 216 46
rect 261 71 263 75
rect 241 62 243 66
rect 251 62 253 66
rect 340 71 342 75
rect 347 71 349 75
rect 357 71 359 75
rect 364 71 366 75
rect 374 71 376 75
rect 397 71 399 75
rect 407 71 409 75
rect 414 71 416 75
rect 424 71 426 75
rect 431 71 433 75
rect 464 71 466 75
rect 474 71 476 75
rect 481 71 483 75
rect 491 71 493 75
rect 498 71 500 75
rect 288 64 290 69
rect 298 64 300 69
rect 308 62 310 66
rect 288 48 290 51
rect 284 46 290 48
rect 284 44 286 46
rect 288 44 290 46
rect 210 42 216 44
rect 177 38 183 40
rect 177 36 179 38
rect 181 36 183 38
rect 112 31 114 33
rect 116 31 121 33
rect 14 17 16 22
rect 24 20 26 25
rect 34 20 36 25
rect 63 16 65 20
rect 112 29 121 31
rect 137 31 139 34
rect 119 26 121 29
rect 129 26 131 30
rect 137 29 141 31
rect 139 26 141 29
rect 146 26 148 35
rect 177 34 183 36
rect 187 38 193 40
rect 187 36 189 38
rect 191 36 193 38
rect 187 34 193 36
rect 177 29 179 34
rect 190 29 192 34
rect 197 29 199 42
rect 214 41 216 42
rect 225 41 227 44
rect 241 41 243 44
rect 214 39 227 41
rect 233 39 243 41
rect 251 40 253 44
rect 261 41 263 44
rect 284 42 290 44
rect 217 31 219 39
rect 233 35 235 39
rect 226 33 235 35
rect 247 38 253 40
rect 247 36 249 38
rect 251 36 253 38
rect 247 34 253 36
rect 257 39 263 41
rect 257 37 259 39
rect 261 37 263 39
rect 257 35 263 37
rect 226 31 228 33
rect 230 31 235 33
rect 103 19 105 22
rect 76 13 78 18
rect 83 13 85 18
rect 103 17 108 19
rect 106 9 108 17
rect 119 13 121 17
rect 129 9 131 17
rect 177 16 179 20
rect 226 29 235 31
rect 251 31 253 34
rect 233 26 235 29
rect 243 26 245 30
rect 251 29 255 31
rect 253 26 255 29
rect 260 26 262 35
rect 288 29 290 42
rect 298 40 300 51
rect 323 58 329 60
rect 323 56 325 58
rect 327 56 329 58
rect 323 54 332 56
rect 330 51 332 54
rect 308 40 310 44
rect 294 38 300 40
rect 294 36 296 38
rect 298 36 300 38
rect 294 34 300 36
rect 304 38 310 40
rect 304 36 306 38
rect 308 36 310 38
rect 304 34 310 36
rect 295 29 297 34
rect 308 29 310 34
rect 217 19 219 22
rect 139 9 141 14
rect 146 9 148 14
rect 106 7 131 9
rect 190 13 192 18
rect 197 13 199 18
rect 217 17 222 19
rect 220 9 222 17
rect 233 13 235 17
rect 243 9 245 17
rect 330 25 332 43
rect 340 40 342 55
rect 347 50 349 55
rect 346 48 352 50
rect 346 46 348 48
rect 350 46 352 48
rect 346 44 352 46
rect 357 40 359 55
rect 364 45 366 55
rect 444 58 450 60
rect 444 56 446 58
rect 448 56 450 58
rect 336 38 342 40
rect 336 36 338 38
rect 340 36 342 38
rect 336 34 342 36
rect 340 25 342 34
rect 347 38 359 40
rect 363 43 369 45
rect 363 41 365 43
rect 367 41 369 43
rect 363 39 369 41
rect 347 25 349 38
rect 353 32 359 34
rect 353 30 355 32
rect 357 30 359 32
rect 353 28 359 30
rect 357 25 359 28
rect 364 25 366 39
rect 374 35 376 53
rect 397 35 399 53
rect 407 45 409 55
rect 404 43 410 45
rect 404 41 406 43
rect 408 41 410 43
rect 404 39 410 41
rect 414 40 416 55
rect 424 50 426 55
rect 421 48 427 50
rect 421 46 423 48
rect 425 46 427 48
rect 421 44 427 46
rect 431 40 433 55
rect 441 54 450 56
rect 441 51 443 54
rect 543 71 545 75
rect 550 71 552 75
rect 572 71 574 75
rect 530 61 532 66
rect 511 58 517 60
rect 511 56 513 58
rect 515 56 517 58
rect 371 33 377 35
rect 371 31 373 33
rect 375 31 377 33
rect 371 29 377 31
rect 396 33 402 35
rect 396 31 398 33
rect 400 31 402 33
rect 396 29 402 31
rect 374 26 376 29
rect 397 26 399 29
rect 253 9 255 14
rect 260 9 262 14
rect 288 13 290 18
rect 295 13 297 18
rect 220 7 245 9
rect 308 16 310 20
rect 330 9 332 19
rect 407 25 409 39
rect 414 38 426 40
rect 414 32 420 34
rect 414 30 416 32
rect 418 30 420 32
rect 414 28 420 30
rect 414 25 416 28
rect 424 25 426 38
rect 431 38 437 40
rect 431 36 433 38
rect 435 36 437 38
rect 431 34 437 36
rect 431 25 433 34
rect 441 25 443 43
rect 464 35 466 53
rect 474 45 476 55
rect 471 43 477 45
rect 471 41 473 43
rect 475 41 477 43
rect 471 39 477 41
rect 481 40 483 55
rect 491 50 493 55
rect 488 48 494 50
rect 488 46 490 48
rect 492 46 494 48
rect 488 44 494 46
rect 498 40 500 55
rect 508 54 517 56
rect 508 51 510 54
rect 463 33 469 35
rect 463 31 465 33
rect 467 31 469 33
rect 463 29 469 31
rect 464 26 466 29
rect 340 13 342 17
rect 347 9 349 17
rect 357 12 359 17
rect 364 12 366 17
rect 374 12 376 17
rect 397 12 399 17
rect 407 12 409 17
rect 414 12 416 17
rect 330 7 349 9
rect 424 9 426 17
rect 431 13 433 17
rect 441 9 443 19
rect 474 25 476 39
rect 481 38 493 40
rect 481 32 487 34
rect 481 30 483 32
rect 485 30 487 32
rect 481 28 487 30
rect 481 25 483 28
rect 491 25 493 38
rect 498 38 504 40
rect 498 36 500 38
rect 502 36 504 38
rect 498 34 504 36
rect 498 25 500 34
rect 508 25 510 43
rect 530 40 532 43
rect 543 40 545 50
rect 550 47 552 50
rect 550 45 556 47
rect 550 43 552 45
rect 554 43 556 45
rect 608 71 610 75
rect 582 62 584 66
rect 592 62 594 66
rect 619 46 625 48
rect 619 44 621 46
rect 623 44 625 46
rect 550 41 556 43
rect 572 41 574 44
rect 530 38 536 40
rect 530 36 532 38
rect 534 36 536 38
rect 530 34 536 36
rect 540 38 546 40
rect 540 36 542 38
rect 544 36 546 38
rect 540 34 546 36
rect 530 31 532 34
rect 540 31 542 34
rect 550 31 552 41
rect 572 39 578 41
rect 572 37 574 39
rect 576 37 578 39
rect 572 35 578 37
rect 582 40 584 44
rect 592 41 594 44
rect 608 41 610 44
rect 619 42 625 44
rect 619 41 621 42
rect 582 38 588 40
rect 592 39 602 41
rect 608 39 621 41
rect 582 36 584 38
rect 586 36 588 38
rect 573 26 575 35
rect 582 34 588 36
rect 600 35 602 39
rect 582 31 584 34
rect 580 29 584 31
rect 600 33 609 35
rect 600 31 605 33
rect 607 31 609 33
rect 616 31 618 39
rect 580 26 582 29
rect 590 26 592 30
rect 600 29 609 31
rect 600 26 602 29
rect 464 12 466 17
rect 474 12 476 17
rect 481 12 483 17
rect 424 7 443 9
rect 491 9 493 17
rect 498 13 500 17
rect 508 9 510 19
rect 530 17 532 22
rect 540 20 542 25
rect 550 20 552 25
rect 491 7 510 9
rect 616 19 618 22
rect 613 17 618 19
rect 573 9 575 14
rect 580 9 582 14
rect 590 9 592 17
rect 600 13 602 17
rect 613 9 615 17
rect 590 7 615 9
<< ndif >>
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 9 22 14 25
rect 16 25 24 31
rect 26 29 34 31
rect 26 27 29 29
rect 31 27 34 29
rect 26 25 34 27
rect 36 25 43 31
rect 96 29 103 31
rect 58 26 63 29
rect 16 22 22 25
rect 18 18 22 22
rect 38 18 43 25
rect 56 24 63 26
rect 56 22 58 24
rect 60 22 63 24
rect 56 20 63 22
rect 65 20 76 29
rect 18 16 24 18
rect 18 14 20 16
rect 22 14 24 16
rect 18 12 24 14
rect 37 16 43 18
rect 67 18 76 20
rect 78 18 83 29
rect 85 24 90 29
rect 96 27 98 29
rect 100 27 103 29
rect 96 25 103 27
rect 85 22 92 24
rect 98 22 103 25
rect 105 26 110 31
rect 210 29 217 31
rect 172 26 177 29
rect 105 22 119 26
rect 85 20 88 22
rect 90 20 92 22
rect 85 18 92 20
rect 110 21 119 22
rect 110 19 112 21
rect 114 19 119 21
rect 37 14 39 16
rect 41 14 43 16
rect 37 12 43 14
rect 67 12 74 18
rect 110 17 119 19
rect 121 24 129 26
rect 121 22 124 24
rect 126 22 129 24
rect 121 17 129 22
rect 131 22 139 26
rect 131 20 134 22
rect 136 20 139 22
rect 131 17 139 20
rect 67 10 69 12
rect 71 10 74 12
rect 67 8 74 10
rect 134 14 139 17
rect 141 14 146 26
rect 148 14 156 26
rect 170 24 177 26
rect 170 22 172 24
rect 174 22 177 24
rect 170 20 177 22
rect 179 20 190 29
rect 181 18 190 20
rect 192 18 197 29
rect 199 24 204 29
rect 210 27 212 29
rect 214 27 217 29
rect 210 25 217 27
rect 199 22 206 24
rect 212 22 217 25
rect 219 26 224 31
rect 219 22 233 26
rect 199 20 202 22
rect 204 20 206 22
rect 199 18 206 20
rect 224 21 233 22
rect 224 19 226 21
rect 228 19 233 21
rect 150 12 156 14
rect 150 10 152 12
rect 154 10 156 12
rect 150 8 156 10
rect 181 12 188 18
rect 224 17 233 19
rect 235 24 243 26
rect 235 22 238 24
rect 240 22 243 24
rect 235 17 243 22
rect 245 22 253 26
rect 245 20 248 22
rect 250 20 253 22
rect 245 17 253 20
rect 181 10 183 12
rect 185 10 188 12
rect 181 8 188 10
rect 248 14 253 17
rect 255 14 260 26
rect 262 14 270 26
rect 283 24 288 29
rect 281 22 288 24
rect 281 20 283 22
rect 285 20 288 22
rect 281 18 288 20
rect 290 18 295 29
rect 297 20 308 29
rect 310 26 315 29
rect 310 24 317 26
rect 369 25 374 26
rect 310 22 313 24
rect 315 22 317 24
rect 310 20 317 22
rect 323 23 330 25
rect 323 21 325 23
rect 327 21 330 23
rect 297 18 306 20
rect 264 12 270 14
rect 264 10 266 12
rect 268 10 270 12
rect 264 8 270 10
rect 299 12 306 18
rect 323 19 330 21
rect 332 23 340 25
rect 332 21 335 23
rect 337 21 340 23
rect 332 19 340 21
rect 299 10 302 12
rect 304 10 306 12
rect 299 8 306 10
rect 334 17 340 19
rect 342 17 347 25
rect 349 21 357 25
rect 349 19 352 21
rect 354 19 357 21
rect 349 17 357 19
rect 359 17 364 25
rect 366 21 374 25
rect 366 19 369 21
rect 371 19 374 21
rect 366 17 374 19
rect 376 24 383 26
rect 376 22 379 24
rect 381 22 383 24
rect 376 20 383 22
rect 390 24 397 26
rect 390 22 392 24
rect 394 22 397 24
rect 390 20 397 22
rect 376 17 381 20
rect 392 17 397 20
rect 399 25 404 26
rect 399 21 407 25
rect 399 19 402 21
rect 404 19 407 21
rect 399 17 407 19
rect 409 17 414 25
rect 416 21 424 25
rect 416 19 419 21
rect 421 19 424 21
rect 416 17 424 19
rect 426 17 431 25
rect 433 23 441 25
rect 433 21 436 23
rect 438 21 441 23
rect 433 19 441 21
rect 443 23 450 25
rect 443 21 446 23
rect 448 21 450 23
rect 443 19 450 21
rect 457 24 464 26
rect 457 22 459 24
rect 461 22 464 24
rect 457 20 464 22
rect 433 17 439 19
rect 459 17 464 20
rect 466 25 471 26
rect 523 29 530 31
rect 523 27 525 29
rect 527 27 530 29
rect 523 25 530 27
rect 466 21 474 25
rect 466 19 469 21
rect 471 19 474 21
rect 466 17 474 19
rect 476 17 481 25
rect 483 21 491 25
rect 483 19 486 21
rect 488 19 491 21
rect 483 17 491 19
rect 493 17 498 25
rect 500 23 508 25
rect 500 21 503 23
rect 505 21 508 23
rect 500 19 508 21
rect 510 23 517 25
rect 510 21 513 23
rect 515 21 517 23
rect 525 22 530 25
rect 532 25 540 31
rect 542 29 550 31
rect 542 27 545 29
rect 547 27 550 29
rect 542 25 550 27
rect 552 25 559 31
rect 611 26 616 31
rect 532 22 538 25
rect 510 19 517 21
rect 500 17 506 19
rect 534 18 538 22
rect 554 18 559 25
rect 534 16 540 18
rect 534 14 536 16
rect 538 14 540 16
rect 534 12 540 14
rect 553 16 559 18
rect 553 14 555 16
rect 557 14 559 16
rect 553 12 559 14
rect 565 14 573 26
rect 575 14 580 26
rect 582 22 590 26
rect 582 20 585 22
rect 587 20 590 22
rect 582 17 590 20
rect 592 24 600 26
rect 592 22 595 24
rect 597 22 600 24
rect 592 17 600 22
rect 602 22 616 26
rect 618 29 625 31
rect 618 27 621 29
rect 623 27 625 29
rect 618 25 625 27
rect 618 22 623 25
rect 602 21 611 22
rect 602 19 607 21
rect 609 19 611 21
rect 602 17 611 19
rect 582 14 587 17
rect 565 12 571 14
rect 565 10 567 12
rect 569 10 571 12
rect 565 8 571 10
<< pdif >>
rect 18 69 27 71
rect 18 67 20 69
rect 22 67 27 69
rect 18 61 27 67
rect 7 59 14 61
rect 7 57 9 59
rect 11 57 14 59
rect 7 52 14 57
rect 7 50 9 52
rect 11 50 14 52
rect 7 48 14 50
rect 9 43 14 48
rect 16 50 27 61
rect 29 50 34 71
rect 36 64 41 71
rect 36 62 43 64
rect 67 62 73 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 58 43 60
rect 36 50 41 58
rect 58 57 63 62
rect 56 55 63 57
rect 56 53 58 55
rect 60 53 63 55
rect 16 43 24 50
rect 56 48 63 53
rect 56 46 58 48
rect 60 46 63 48
rect 56 44 63 46
rect 65 60 73 62
rect 65 58 68 60
rect 70 58 73 60
rect 65 51 73 58
rect 75 62 83 64
rect 75 60 78 62
rect 80 60 83 62
rect 75 55 83 60
rect 75 53 78 55
rect 80 53 83 55
rect 75 51 83 53
rect 85 62 92 64
rect 85 60 88 62
rect 90 60 92 62
rect 85 51 92 60
rect 65 44 71 51
rect 106 50 111 71
rect 104 48 111 50
rect 104 46 106 48
rect 108 46 111 48
rect 104 44 111 46
rect 113 69 125 71
rect 113 67 116 69
rect 118 67 125 69
rect 113 62 125 67
rect 142 62 147 71
rect 113 60 116 62
rect 118 60 127 62
rect 113 44 127 60
rect 129 55 137 62
rect 129 53 132 55
rect 134 53 137 55
rect 129 48 137 53
rect 129 46 132 48
rect 134 46 137 48
rect 129 44 137 46
rect 139 55 147 62
rect 139 53 142 55
rect 144 53 147 55
rect 139 44 147 53
rect 149 65 154 71
rect 149 63 156 65
rect 149 61 152 63
rect 154 61 156 63
rect 181 62 187 64
rect 149 59 156 61
rect 149 44 154 59
rect 172 57 177 62
rect 170 55 177 57
rect 170 53 172 55
rect 174 53 177 55
rect 170 48 177 53
rect 170 46 172 48
rect 174 46 177 48
rect 170 44 177 46
rect 179 60 187 62
rect 179 58 182 60
rect 184 58 187 60
rect 179 51 187 58
rect 189 62 197 64
rect 189 60 192 62
rect 194 60 197 62
rect 189 55 197 60
rect 189 53 192 55
rect 194 53 197 55
rect 189 51 197 53
rect 199 62 206 64
rect 199 60 202 62
rect 204 60 206 62
rect 199 51 206 60
rect 179 44 185 51
rect 220 50 225 71
rect 218 48 225 50
rect 218 46 220 48
rect 222 46 225 48
rect 218 44 225 46
rect 227 69 239 71
rect 227 67 230 69
rect 232 67 239 69
rect 227 62 239 67
rect 256 62 261 71
rect 227 60 230 62
rect 232 60 241 62
rect 227 44 241 60
rect 243 55 251 62
rect 243 53 246 55
rect 248 53 251 55
rect 243 48 251 53
rect 243 46 246 48
rect 248 46 251 48
rect 243 44 251 46
rect 253 55 261 62
rect 253 53 256 55
rect 258 53 261 55
rect 253 44 261 53
rect 263 65 268 71
rect 263 63 270 65
rect 333 69 340 71
rect 333 67 335 69
rect 337 67 340 69
rect 263 61 266 63
rect 268 61 270 63
rect 263 59 270 61
rect 281 62 288 64
rect 281 60 283 62
rect 285 60 288 62
rect 263 44 268 59
rect 281 51 288 60
rect 290 62 298 64
rect 290 60 293 62
rect 295 60 298 62
rect 290 55 298 60
rect 290 53 293 55
rect 295 53 298 55
rect 290 51 298 53
rect 300 62 306 64
rect 300 60 308 62
rect 300 58 303 60
rect 305 58 308 60
rect 300 51 308 58
rect 302 44 308 51
rect 310 57 315 62
rect 333 59 340 67
rect 310 55 317 57
rect 310 53 313 55
rect 315 53 317 55
rect 310 48 317 53
rect 334 55 340 59
rect 342 55 347 71
rect 349 59 357 71
rect 349 57 352 59
rect 354 57 357 59
rect 349 55 357 57
rect 359 55 364 71
rect 366 69 374 71
rect 366 67 369 69
rect 371 67 374 69
rect 366 55 374 67
rect 334 51 338 55
rect 325 49 330 51
rect 310 46 313 48
rect 315 46 317 48
rect 310 44 317 46
rect 323 47 330 49
rect 323 45 325 47
rect 327 45 330 47
rect 323 43 330 45
rect 332 43 338 51
rect 369 53 374 55
rect 376 64 381 71
rect 392 64 397 71
rect 376 62 383 64
rect 376 60 379 62
rect 381 60 383 62
rect 376 58 383 60
rect 390 62 397 64
rect 390 60 392 62
rect 394 60 397 62
rect 390 58 397 60
rect 376 53 381 58
rect 392 53 397 58
rect 399 69 407 71
rect 399 67 402 69
rect 404 67 407 69
rect 399 55 407 67
rect 409 55 414 71
rect 416 59 424 71
rect 416 57 419 59
rect 421 57 424 59
rect 416 55 424 57
rect 426 55 431 71
rect 433 69 440 71
rect 433 67 436 69
rect 438 67 440 69
rect 433 59 440 67
rect 459 64 464 71
rect 457 62 464 64
rect 457 60 459 62
rect 461 60 464 62
rect 433 55 439 59
rect 457 58 464 60
rect 399 53 404 55
rect 435 51 439 55
rect 459 53 464 58
rect 466 69 474 71
rect 466 67 469 69
rect 471 67 474 69
rect 466 55 474 67
rect 476 55 481 71
rect 483 59 491 71
rect 483 57 486 59
rect 488 57 491 59
rect 483 55 491 57
rect 493 55 498 71
rect 500 69 507 71
rect 500 67 503 69
rect 505 67 507 69
rect 534 69 543 71
rect 500 59 507 67
rect 534 67 536 69
rect 538 67 543 69
rect 534 61 543 67
rect 500 55 506 59
rect 466 53 471 55
rect 435 43 441 51
rect 443 49 448 51
rect 443 47 450 49
rect 443 45 446 47
rect 448 45 450 47
rect 443 43 450 45
rect 502 51 506 55
rect 523 59 530 61
rect 523 57 525 59
rect 527 57 530 59
rect 523 52 530 57
rect 502 43 508 51
rect 510 49 515 51
rect 523 50 525 52
rect 527 50 530 52
rect 510 47 517 49
rect 523 48 530 50
rect 510 45 513 47
rect 515 45 517 47
rect 510 43 517 45
rect 525 43 530 48
rect 532 50 543 61
rect 545 50 550 71
rect 552 64 557 71
rect 567 65 572 71
rect 552 62 559 64
rect 552 60 555 62
rect 557 60 559 62
rect 552 58 559 60
rect 565 63 572 65
rect 565 61 567 63
rect 569 61 572 63
rect 565 59 572 61
rect 552 50 557 58
rect 532 43 540 50
rect 567 44 572 59
rect 574 62 579 71
rect 596 69 608 71
rect 596 67 603 69
rect 605 67 608 69
rect 596 62 608 67
rect 574 55 582 62
rect 574 53 577 55
rect 579 53 582 55
rect 574 44 582 53
rect 584 55 592 62
rect 584 53 587 55
rect 589 53 592 55
rect 584 48 592 53
rect 584 46 587 48
rect 589 46 592 48
rect 584 44 592 46
rect 594 60 603 62
rect 605 60 608 62
rect 594 44 608 60
rect 610 50 615 71
rect 610 48 617 50
rect 610 46 613 48
rect 615 46 617 48
rect 610 44 617 46
<< alu1 >>
rect 3 72 633 77
rect 3 70 10 72
rect 12 70 59 72
rect 61 70 132 72
rect 134 70 173 72
rect 175 70 246 72
rect 248 70 312 72
rect 314 70 526 72
rect 528 70 587 72
rect 589 70 633 72
rect 3 69 633 70
rect 7 63 11 64
rect 7 59 20 63
rect 7 57 9 59
rect 7 52 11 57
rect 7 50 9 52
rect 7 31 11 50
rect 39 53 43 56
rect 56 55 61 57
rect 56 53 58 55
rect 60 53 61 55
rect 96 58 108 64
rect 39 49 61 53
rect 39 47 43 49
rect 22 45 43 47
rect 22 43 36 45
rect 38 43 43 45
rect 56 48 61 49
rect 56 46 58 48
rect 60 46 61 48
rect 56 44 61 46
rect 88 53 92 56
rect 88 51 89 53
rect 91 51 92 53
rect 7 29 12 31
rect 7 27 9 29
rect 11 27 12 29
rect 7 25 12 27
rect 22 38 43 39
rect 22 36 26 38
rect 28 36 40 38
rect 42 36 43 38
rect 22 35 43 36
rect 39 26 43 35
rect 56 24 60 44
rect 88 47 92 51
rect 79 46 92 47
rect 79 44 85 46
rect 87 44 92 46
rect 79 43 92 44
rect 96 53 101 58
rect 96 51 98 53
rect 100 51 101 53
rect 96 46 101 51
rect 96 44 98 46
rect 100 44 101 46
rect 96 42 101 44
rect 71 38 85 39
rect 71 36 75 38
rect 77 36 85 38
rect 71 35 85 36
rect 56 22 58 24
rect 60 22 68 24
rect 56 18 68 22
rect 80 29 85 35
rect 80 27 81 29
rect 83 27 85 29
rect 80 26 85 27
rect 112 33 117 40
rect 140 55 156 56
rect 140 53 142 55
rect 144 53 156 55
rect 140 51 156 53
rect 112 32 114 33
rect 104 31 114 32
rect 116 31 117 33
rect 104 29 117 31
rect 104 27 106 29
rect 108 27 117 29
rect 104 26 117 27
rect 152 30 156 51
rect 152 28 153 30
rect 155 28 156 30
rect 152 23 156 28
rect 132 22 156 23
rect 132 20 134 22
rect 136 20 156 22
rect 132 19 156 20
rect 170 55 175 57
rect 170 53 172 55
rect 174 53 175 55
rect 210 58 222 64
rect 170 48 175 53
rect 170 46 172 48
rect 174 46 175 48
rect 170 44 175 46
rect 202 53 206 56
rect 202 51 203 53
rect 205 51 206 53
rect 170 38 174 44
rect 170 36 171 38
rect 173 36 174 38
rect 170 24 174 36
rect 202 47 206 51
rect 193 46 206 47
rect 193 44 199 46
rect 201 44 206 46
rect 193 43 206 44
rect 210 53 215 58
rect 210 51 212 53
rect 214 51 215 53
rect 210 46 215 51
rect 210 44 212 46
rect 214 44 215 46
rect 210 42 215 44
rect 185 38 199 39
rect 185 36 189 38
rect 191 36 199 38
rect 185 35 199 36
rect 170 22 172 24
rect 174 22 182 24
rect 170 18 182 22
rect 194 29 199 35
rect 194 27 195 29
rect 197 27 199 29
rect 194 26 199 27
rect 226 33 231 40
rect 254 55 270 56
rect 254 53 256 55
rect 258 53 270 55
rect 254 51 270 53
rect 266 45 270 51
rect 266 43 267 45
rect 269 43 270 45
rect 281 47 285 56
rect 323 58 328 64
rect 370 62 383 63
rect 370 60 379 62
rect 381 60 383 62
rect 312 55 317 57
rect 281 46 294 47
rect 281 44 286 46
rect 288 44 294 46
rect 281 43 294 44
rect 226 32 228 33
rect 218 31 228 32
rect 230 31 231 33
rect 218 29 231 31
rect 218 27 220 29
rect 222 27 231 29
rect 218 26 231 27
rect 266 23 270 43
rect 288 38 302 39
rect 288 36 296 38
rect 298 36 302 38
rect 288 35 302 36
rect 312 53 313 55
rect 315 53 317 55
rect 312 48 317 53
rect 323 56 325 58
rect 327 56 328 58
rect 370 59 383 60
rect 323 55 328 56
rect 323 54 336 55
rect 323 52 333 54
rect 335 52 336 54
rect 323 51 336 52
rect 312 46 313 48
rect 315 46 317 48
rect 312 44 317 46
rect 288 26 293 35
rect 313 30 317 44
rect 313 28 314 30
rect 316 28 317 30
rect 313 24 317 28
rect 246 22 270 23
rect 246 20 248 22
rect 250 20 270 22
rect 246 19 270 20
rect 305 22 313 24
rect 315 22 317 24
rect 305 18 317 22
rect 337 38 343 40
rect 337 36 338 38
rect 340 36 343 38
rect 337 31 343 36
rect 330 30 343 31
rect 330 28 331 30
rect 333 28 343 30
rect 355 46 367 48
rect 355 44 356 46
rect 358 44 367 46
rect 355 43 367 44
rect 355 42 365 43
rect 363 41 365 42
rect 363 34 367 41
rect 379 38 383 59
rect 379 36 380 38
rect 382 36 383 38
rect 330 27 343 28
rect 379 26 383 36
rect 378 24 383 26
rect 378 22 379 24
rect 381 22 383 24
rect 378 20 383 22
rect 379 18 383 20
rect 390 62 403 63
rect 390 60 392 62
rect 394 60 403 62
rect 390 59 403 60
rect 390 26 394 59
rect 445 58 450 64
rect 445 56 446 58
rect 448 56 450 58
rect 445 55 450 56
rect 437 51 450 55
rect 457 62 470 63
rect 457 60 459 62
rect 461 60 470 62
rect 457 59 470 60
rect 406 43 418 48
rect 408 42 418 43
rect 408 41 410 42
rect 406 38 410 41
rect 406 36 407 38
rect 409 36 410 38
rect 406 34 410 36
rect 430 38 436 40
rect 430 36 433 38
rect 435 36 436 38
rect 430 31 436 36
rect 430 30 443 31
rect 430 28 438 30
rect 440 28 443 30
rect 430 27 443 28
rect 390 24 395 26
rect 390 22 392 24
rect 394 22 395 24
rect 390 20 395 22
rect 390 18 394 20
rect 457 30 461 59
rect 512 58 517 64
rect 512 56 513 58
rect 515 56 517 58
rect 512 55 517 56
rect 504 54 517 55
rect 504 52 505 54
rect 507 52 517 54
rect 504 51 517 52
rect 523 63 527 64
rect 523 59 536 63
rect 523 57 525 59
rect 523 52 527 57
rect 523 50 525 52
rect 473 45 485 48
rect 473 43 481 45
rect 483 43 485 45
rect 475 42 485 43
rect 475 41 477 42
rect 457 28 458 30
rect 460 28 461 30
rect 473 34 477 41
rect 457 26 461 28
rect 497 38 503 40
rect 497 36 500 38
rect 502 36 503 38
rect 497 31 503 36
rect 497 30 510 31
rect 497 28 506 30
rect 508 28 510 30
rect 497 27 510 28
rect 457 24 462 26
rect 457 22 459 24
rect 461 22 462 24
rect 457 20 462 22
rect 457 18 461 20
rect 523 46 527 50
rect 523 44 524 46
rect 526 44 527 46
rect 523 31 527 44
rect 555 47 559 56
rect 538 45 559 47
rect 538 43 552 45
rect 554 43 559 45
rect 565 55 581 56
rect 565 53 577 55
rect 579 53 581 55
rect 565 51 581 53
rect 523 29 528 31
rect 523 27 525 29
rect 527 27 528 29
rect 523 25 528 27
rect 538 38 559 39
rect 538 36 542 38
rect 544 36 559 38
rect 538 35 559 36
rect 555 26 559 35
rect 565 30 569 51
rect 613 58 625 64
rect 565 28 566 30
rect 568 28 569 30
rect 565 23 569 28
rect 604 33 609 40
rect 620 46 625 58
rect 620 44 621 46
rect 623 44 625 46
rect 620 42 625 44
rect 604 31 605 33
rect 607 32 609 33
rect 607 31 617 32
rect 604 26 617 31
rect 565 22 589 23
rect 565 20 585 22
rect 587 20 589 22
rect 565 19 589 20
rect 3 12 633 13
rect 3 10 10 12
rect 12 10 59 12
rect 61 10 69 12
rect 71 10 99 12
rect 101 10 152 12
rect 154 10 173 12
rect 175 10 183 12
rect 185 10 213 12
rect 215 10 266 12
rect 268 10 302 12
rect 304 10 312 12
rect 314 10 526 12
rect 528 10 567 12
rect 569 10 620 12
rect 622 10 633 12
rect 3 5 633 10
<< alu2 >>
rect 332 54 509 55
rect 88 53 101 54
rect 88 51 89 53
rect 91 51 98 53
rect 100 51 101 53
rect 88 50 101 51
rect 202 53 215 54
rect 202 51 203 53
rect 205 51 212 53
rect 214 51 215 53
rect 332 52 333 54
rect 335 52 505 54
rect 507 52 509 54
rect 332 51 509 52
rect 202 50 215 51
rect 266 46 360 47
rect 266 45 356 46
rect 266 43 267 45
rect 269 44 356 45
rect 358 44 360 46
rect 269 43 360 44
rect 266 42 360 43
rect 480 46 527 47
rect 480 45 524 46
rect 480 43 481 45
rect 483 44 524 45
rect 526 44 527 46
rect 483 43 527 44
rect 480 42 527 43
rect 39 38 174 39
rect 39 36 40 38
rect 42 36 171 38
rect 173 36 174 38
rect 39 35 174 36
rect 379 38 410 39
rect 379 36 380 38
rect 382 36 407 38
rect 409 36 410 38
rect 379 35 410 36
rect 80 29 112 31
rect 80 27 81 29
rect 83 27 106 29
rect 108 27 112 29
rect 80 26 112 27
rect 152 30 226 31
rect 152 28 153 30
rect 155 29 226 30
rect 155 28 195 29
rect 152 27 195 28
rect 197 27 220 29
rect 222 27 226 29
rect 313 30 334 31
rect 313 28 314 30
rect 316 28 331 30
rect 333 28 334 30
rect 313 27 334 28
rect 437 30 461 31
rect 437 28 438 30
rect 440 28 458 30
rect 460 28 461 30
rect 437 27 461 28
rect 505 30 569 31
rect 505 28 506 30
rect 508 28 566 30
rect 568 28 569 30
rect 505 27 569 28
rect 152 26 226 27
<< ptie >>
rect 8 12 14 14
rect 57 12 63 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 57 10 59 12
rect 61 10 63 12
rect 57 8 63 10
rect 97 12 103 14
rect 97 10 99 12
rect 101 10 103 12
rect 97 8 103 10
rect 171 12 177 14
rect 171 10 173 12
rect 175 10 177 12
rect 171 8 177 10
rect 211 12 217 14
rect 211 10 213 12
rect 215 10 217 12
rect 211 8 217 10
rect 310 12 316 14
rect 310 10 312 12
rect 314 10 316 12
rect 310 8 316 10
rect 524 12 530 14
rect 524 10 526 12
rect 528 10 530 12
rect 524 8 530 10
rect 618 12 624 14
rect 618 10 620 12
rect 622 10 624 12
rect 618 8 624 10
<< ntie >>
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 57 72 63 74
rect 8 68 14 70
rect 57 70 59 72
rect 61 70 63 72
rect 130 72 136 74
rect 57 68 63 70
rect 130 70 132 72
rect 134 70 136 72
rect 171 72 177 74
rect 130 68 136 70
rect 171 70 173 72
rect 175 70 177 72
rect 244 72 250 74
rect 171 68 177 70
rect 244 70 246 72
rect 248 70 250 72
rect 310 72 316 74
rect 244 68 250 70
rect 310 70 312 72
rect 314 70 316 72
rect 524 72 530 74
rect 310 68 316 70
rect 524 70 526 72
rect 528 70 530 72
rect 585 72 591 74
rect 524 68 530 70
rect 585 70 587 72
rect 589 70 591 72
rect 585 68 591 70
<< nmos >>
rect 14 22 16 31
rect 24 25 26 31
rect 34 25 36 31
rect 63 20 65 29
rect 76 18 78 29
rect 83 18 85 29
rect 103 22 105 31
rect 119 17 121 26
rect 129 17 131 26
rect 139 14 141 26
rect 146 14 148 26
rect 177 20 179 29
rect 190 18 192 29
rect 197 18 199 29
rect 217 22 219 31
rect 233 17 235 26
rect 243 17 245 26
rect 253 14 255 26
rect 260 14 262 26
rect 288 18 290 29
rect 295 18 297 29
rect 308 20 310 29
rect 330 19 332 25
rect 340 17 342 25
rect 347 17 349 25
rect 357 17 359 25
rect 364 17 366 25
rect 374 17 376 26
rect 397 17 399 26
rect 407 17 409 25
rect 414 17 416 25
rect 424 17 426 25
rect 431 17 433 25
rect 441 19 443 25
rect 464 17 466 26
rect 474 17 476 25
rect 481 17 483 25
rect 491 17 493 25
rect 498 17 500 25
rect 508 19 510 25
rect 530 22 532 31
rect 540 25 542 31
rect 550 25 552 31
rect 573 14 575 26
rect 580 14 582 26
rect 590 17 592 26
rect 600 17 602 26
rect 616 22 618 31
<< pmos >>
rect 14 43 16 61
rect 27 50 29 71
rect 34 50 36 71
rect 63 44 65 62
rect 73 51 75 64
rect 83 51 85 64
rect 111 44 113 71
rect 127 44 129 62
rect 137 44 139 62
rect 147 44 149 71
rect 177 44 179 62
rect 187 51 189 64
rect 197 51 199 64
rect 225 44 227 71
rect 241 44 243 62
rect 251 44 253 62
rect 261 44 263 71
rect 288 51 290 64
rect 298 51 300 64
rect 308 44 310 62
rect 340 55 342 71
rect 347 55 349 71
rect 357 55 359 71
rect 364 55 366 71
rect 330 43 332 51
rect 374 53 376 71
rect 397 53 399 71
rect 407 55 409 71
rect 414 55 416 71
rect 424 55 426 71
rect 431 55 433 71
rect 464 53 466 71
rect 474 55 476 71
rect 481 55 483 71
rect 491 55 493 71
rect 498 55 500 71
rect 441 43 443 51
rect 508 43 510 51
rect 530 43 532 61
rect 543 50 545 71
rect 550 50 552 71
rect 572 44 574 71
rect 582 44 584 62
rect 592 44 594 62
rect 608 44 610 71
<< polyct0 >>
rect 16 36 18 38
rect 65 36 67 38
rect 135 36 137 38
rect 145 37 147 39
rect 179 36 181 38
rect 249 36 251 38
rect 259 37 261 39
rect 306 36 308 38
rect 348 46 350 48
rect 355 30 357 32
rect 423 46 425 48
rect 373 31 375 33
rect 398 31 400 33
rect 416 30 418 32
rect 490 46 492 48
rect 465 31 467 33
rect 483 30 485 32
rect 532 36 534 38
rect 574 37 576 39
rect 584 36 586 38
<< polyct1 >>
rect 36 43 38 45
rect 26 36 28 38
rect 85 44 87 46
rect 98 44 100 46
rect 75 36 77 38
rect 199 44 201 46
rect 212 44 214 46
rect 286 44 288 46
rect 114 31 116 33
rect 189 36 191 38
rect 228 31 230 33
rect 325 56 327 58
rect 296 36 298 38
rect 446 56 448 58
rect 338 36 340 38
rect 365 41 367 43
rect 406 41 408 43
rect 513 56 515 58
rect 433 36 435 38
rect 473 41 475 43
rect 500 36 502 38
rect 552 43 554 45
rect 621 44 623 46
rect 542 36 544 38
rect 605 31 607 33
<< ndifct0 >>
rect 29 27 31 29
rect 20 14 22 16
rect 98 27 100 29
rect 88 20 90 22
rect 112 19 114 21
rect 39 14 41 16
rect 124 22 126 24
rect 212 27 214 29
rect 202 20 204 22
rect 226 19 228 21
rect 238 22 240 24
rect 283 20 285 22
rect 325 21 327 23
rect 335 21 337 23
rect 352 19 354 21
rect 369 19 371 21
rect 402 19 404 21
rect 419 19 421 21
rect 436 21 438 23
rect 446 21 448 23
rect 469 19 471 21
rect 486 19 488 21
rect 503 21 505 23
rect 513 21 515 23
rect 545 27 547 29
rect 536 14 538 16
rect 555 14 557 16
rect 595 22 597 24
rect 621 27 623 29
rect 607 19 609 21
<< ndifct1 >>
rect 9 27 11 29
rect 58 22 60 24
rect 134 20 136 22
rect 69 10 71 12
rect 172 22 174 24
rect 152 10 154 12
rect 248 20 250 22
rect 183 10 185 12
rect 313 22 315 24
rect 266 10 268 12
rect 302 10 304 12
rect 379 22 381 24
rect 392 22 394 24
rect 459 22 461 24
rect 525 27 527 29
rect 585 20 587 22
rect 567 10 569 12
<< ntiect1 >>
rect 10 70 12 72
rect 59 70 61 72
rect 132 70 134 72
rect 173 70 175 72
rect 246 70 248 72
rect 312 70 314 72
rect 526 70 528 72
rect 587 70 589 72
<< ptiect1 >>
rect 10 10 12 12
rect 59 10 61 12
rect 99 10 101 12
rect 173 10 175 12
rect 213 10 215 12
rect 312 10 314 12
rect 526 10 528 12
rect 620 10 622 12
<< pdifct0 >>
rect 20 67 22 69
rect 39 60 41 62
rect 68 58 70 60
rect 78 60 80 62
rect 78 53 80 55
rect 88 60 90 62
rect 106 46 108 48
rect 116 67 118 69
rect 116 60 118 62
rect 132 53 134 55
rect 132 46 134 48
rect 152 61 154 63
rect 182 58 184 60
rect 192 60 194 62
rect 192 53 194 55
rect 202 60 204 62
rect 220 46 222 48
rect 230 67 232 69
rect 230 60 232 62
rect 246 53 248 55
rect 246 46 248 48
rect 335 67 337 69
rect 266 61 268 63
rect 283 60 285 62
rect 293 60 295 62
rect 293 53 295 55
rect 303 58 305 60
rect 352 57 354 59
rect 369 67 371 69
rect 325 45 327 47
rect 402 67 404 69
rect 419 57 421 59
rect 436 67 438 69
rect 469 67 471 69
rect 486 57 488 59
rect 503 67 505 69
rect 536 67 538 69
rect 446 45 448 47
rect 513 45 515 47
rect 555 60 557 62
rect 567 61 569 63
rect 603 67 605 69
rect 587 53 589 55
rect 587 46 589 48
rect 603 60 605 62
rect 613 46 615 48
<< pdifct1 >>
rect 9 57 11 59
rect 9 50 11 52
rect 58 53 60 55
rect 58 46 60 48
rect 142 53 144 55
rect 172 53 174 55
rect 172 46 174 48
rect 256 53 258 55
rect 313 53 315 55
rect 313 46 315 48
rect 379 60 381 62
rect 392 60 394 62
rect 459 60 461 62
rect 525 57 527 59
rect 525 50 527 52
rect 577 53 579 55
<< alu0 >>
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 26 62 43 63
rect 26 60 39 62
rect 41 60 43 62
rect 26 59 43 60
rect 66 60 72 69
rect 11 48 12 59
rect 26 55 30 59
rect 66 58 68 60
rect 70 58 72 60
rect 66 57 72 58
rect 77 62 81 64
rect 77 60 78 62
rect 80 60 81 62
rect 15 51 30 55
rect 77 55 81 60
rect 86 62 92 69
rect 115 67 116 69
rect 118 67 119 69
rect 86 60 88 62
rect 90 60 92 62
rect 86 59 92 60
rect 115 62 119 67
rect 115 60 116 62
rect 118 60 119 62
rect 115 58 119 60
rect 123 63 156 64
rect 123 61 152 63
rect 154 61 156 63
rect 123 60 156 61
rect 180 60 186 69
rect 77 54 78 55
rect 15 38 19 51
rect 64 53 78 54
rect 80 53 81 55
rect 64 50 81 53
rect 34 42 40 43
rect 15 36 16 38
rect 18 36 19 38
rect 15 30 19 36
rect 15 29 33 30
rect 15 27 29 29
rect 31 27 33 29
rect 15 26 33 27
rect 64 38 68 50
rect 123 49 127 60
rect 180 58 182 60
rect 184 58 186 60
rect 180 57 186 58
rect 191 62 195 64
rect 191 60 192 62
rect 194 60 195 62
rect 104 48 127 49
rect 104 46 106 48
rect 108 46 127 48
rect 104 45 127 46
rect 104 39 108 45
rect 64 36 65 38
rect 67 36 68 38
rect 64 31 68 36
rect 64 27 76 31
rect 60 24 61 26
rect 72 23 76 27
rect 97 35 108 39
rect 97 29 101 35
rect 123 39 127 45
rect 131 55 135 57
rect 131 53 132 55
rect 134 53 135 55
rect 131 48 135 53
rect 131 46 132 48
rect 134 47 135 48
rect 134 46 147 47
rect 131 43 147 46
rect 143 41 147 43
rect 143 39 148 41
rect 123 38 139 39
rect 123 36 135 38
rect 137 36 139 38
rect 123 35 139 36
rect 143 37 145 39
rect 147 37 148 39
rect 143 35 148 37
rect 97 27 98 29
rect 100 27 101 29
rect 97 25 101 27
rect 143 31 147 35
rect 123 27 147 31
rect 123 24 127 27
rect 72 22 92 23
rect 123 22 124 24
rect 126 22 127 24
rect 72 20 88 22
rect 90 20 92 22
rect 72 19 92 20
rect 110 21 116 22
rect 110 19 112 21
rect 114 19 116 21
rect 123 20 127 22
rect 191 55 195 60
rect 200 62 206 69
rect 229 67 230 69
rect 232 67 233 69
rect 200 60 202 62
rect 204 60 206 62
rect 200 59 206 60
rect 229 62 233 67
rect 229 60 230 62
rect 232 60 233 62
rect 229 58 233 60
rect 237 63 270 64
rect 237 61 266 63
rect 268 61 270 63
rect 237 60 270 61
rect 281 62 287 69
rect 281 60 283 62
rect 285 60 287 62
rect 191 54 192 55
rect 178 53 192 54
rect 194 53 195 55
rect 178 50 195 53
rect 178 38 182 50
rect 237 49 241 60
rect 281 59 287 60
rect 292 62 296 64
rect 292 60 293 62
rect 295 60 296 62
rect 218 48 241 49
rect 218 46 220 48
rect 222 46 241 48
rect 218 45 241 46
rect 218 39 222 45
rect 178 36 179 38
rect 181 36 182 38
rect 178 31 182 36
rect 178 27 190 31
rect 174 24 175 26
rect 18 16 24 17
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 37 16 43 17
rect 37 14 39 16
rect 41 14 43 16
rect 37 13 43 14
rect 110 13 116 19
rect 186 23 190 27
rect 211 35 222 39
rect 211 29 215 35
rect 237 39 241 45
rect 245 55 249 57
rect 245 53 246 55
rect 248 53 249 55
rect 245 48 249 53
rect 245 46 246 48
rect 248 47 249 48
rect 248 46 261 47
rect 245 43 261 46
rect 257 41 261 43
rect 292 55 296 60
rect 301 60 307 69
rect 334 67 335 69
rect 337 67 338 69
rect 334 65 338 67
rect 367 67 369 69
rect 371 67 373 69
rect 367 66 373 67
rect 400 67 402 69
rect 404 67 406 69
rect 400 66 406 67
rect 435 67 436 69
rect 438 67 439 69
rect 435 65 439 67
rect 467 67 469 69
rect 471 67 473 69
rect 467 66 473 67
rect 502 67 503 69
rect 505 67 506 69
rect 502 65 506 67
rect 534 67 536 69
rect 538 67 540 69
rect 534 66 540 67
rect 602 67 603 69
rect 605 67 606 69
rect 301 58 303 60
rect 305 58 307 60
rect 301 57 307 58
rect 292 53 293 55
rect 295 54 296 55
rect 295 53 309 54
rect 292 50 309 53
rect 257 39 262 41
rect 237 38 253 39
rect 237 36 249 38
rect 251 36 253 38
rect 237 35 253 36
rect 257 37 259 39
rect 261 37 262 39
rect 257 35 262 37
rect 211 27 212 29
rect 214 27 215 29
rect 211 25 215 27
rect 257 31 261 35
rect 237 27 261 31
rect 237 24 241 27
rect 186 22 206 23
rect 237 22 238 24
rect 240 22 241 24
rect 305 38 309 50
rect 350 59 363 60
rect 350 57 352 59
rect 354 57 363 59
rect 350 56 363 57
rect 359 52 375 56
rect 347 48 351 50
rect 305 36 306 38
rect 308 36 309 38
rect 305 31 309 36
rect 297 27 309 31
rect 297 23 301 27
rect 312 24 313 26
rect 186 20 202 22
rect 204 20 206 22
rect 186 19 206 20
rect 224 21 230 22
rect 224 19 226 21
rect 228 19 230 21
rect 237 20 241 22
rect 281 22 301 23
rect 281 20 283 22
rect 285 20 301 22
rect 281 19 301 20
rect 224 13 230 19
rect 323 47 348 48
rect 323 45 325 47
rect 327 46 348 47
rect 350 46 351 48
rect 327 45 351 46
rect 323 44 351 45
rect 323 24 327 44
rect 347 34 351 44
rect 367 39 368 45
rect 371 35 375 52
rect 347 32 358 34
rect 347 30 355 32
rect 357 30 358 32
rect 371 33 376 35
rect 371 31 373 33
rect 375 31 376 33
rect 347 28 358 30
rect 361 29 376 31
rect 361 27 375 29
rect 323 23 329 24
rect 323 21 325 23
rect 327 21 329 23
rect 323 20 329 21
rect 333 23 339 24
rect 333 21 335 23
rect 337 21 339 23
rect 361 22 365 27
rect 333 13 339 21
rect 350 21 365 22
rect 350 19 352 21
rect 354 19 365 21
rect 350 18 365 19
rect 368 21 372 23
rect 368 19 369 21
rect 371 19 372 21
rect 368 13 372 19
rect 410 59 423 60
rect 410 57 419 59
rect 421 57 423 59
rect 410 56 423 57
rect 398 52 414 56
rect 398 35 402 52
rect 477 59 490 60
rect 422 48 426 50
rect 405 39 406 45
rect 422 46 423 48
rect 425 47 450 48
rect 425 46 446 47
rect 422 45 446 46
rect 448 45 450 47
rect 422 44 450 45
rect 397 33 402 35
rect 422 34 426 44
rect 397 31 398 33
rect 400 31 402 33
rect 415 32 426 34
rect 397 29 412 31
rect 398 27 412 29
rect 415 30 416 32
rect 418 30 426 32
rect 415 28 426 30
rect 401 21 405 23
rect 401 19 402 21
rect 404 19 405 21
rect 401 13 405 19
rect 408 22 412 27
rect 446 24 450 44
rect 434 23 440 24
rect 408 21 423 22
rect 408 19 419 21
rect 421 19 423 21
rect 408 18 423 19
rect 434 21 436 23
rect 438 21 440 23
rect 434 13 440 21
rect 444 23 450 24
rect 444 21 446 23
rect 448 21 450 23
rect 444 20 450 21
rect 477 57 486 59
rect 488 57 490 59
rect 477 56 490 57
rect 465 52 481 56
rect 465 35 469 52
rect 565 63 598 64
rect 542 62 559 63
rect 542 60 555 62
rect 557 60 559 62
rect 565 61 567 63
rect 569 61 598 63
rect 565 60 598 61
rect 542 59 559 60
rect 489 48 493 50
rect 472 39 473 45
rect 489 46 490 48
rect 492 47 517 48
rect 492 46 513 47
rect 489 45 513 46
rect 515 45 517 47
rect 489 44 517 45
rect 464 33 469 35
rect 489 34 493 44
rect 464 31 465 33
rect 467 31 469 33
rect 482 32 493 34
rect 464 29 479 31
rect 465 27 479 29
rect 482 30 483 32
rect 485 30 493 32
rect 482 28 493 30
rect 468 21 472 23
rect 468 19 469 21
rect 471 19 472 21
rect 468 13 472 19
rect 475 22 479 27
rect 513 24 517 44
rect 527 48 528 59
rect 542 55 546 59
rect 531 51 546 55
rect 531 38 535 51
rect 586 55 590 57
rect 586 53 587 55
rect 589 53 590 55
rect 550 42 556 43
rect 531 36 532 38
rect 534 36 535 38
rect 531 30 535 36
rect 531 29 549 30
rect 531 27 545 29
rect 547 27 549 29
rect 531 26 549 27
rect 586 48 590 53
rect 586 47 587 48
rect 574 46 587 47
rect 589 46 590 48
rect 574 43 590 46
rect 594 49 598 60
rect 602 62 606 67
rect 602 60 603 62
rect 605 60 606 62
rect 602 58 606 60
rect 594 48 617 49
rect 594 46 613 48
rect 615 46 617 48
rect 594 45 617 46
rect 574 41 578 43
rect 573 39 578 41
rect 594 39 598 45
rect 573 37 574 39
rect 576 37 578 39
rect 573 35 578 37
rect 582 38 598 39
rect 582 36 584 38
rect 586 36 598 38
rect 582 35 598 36
rect 501 23 507 24
rect 475 21 490 22
rect 475 19 486 21
rect 488 19 490 21
rect 475 18 490 19
rect 501 21 503 23
rect 505 21 507 23
rect 501 13 507 21
rect 511 23 517 24
rect 511 21 513 23
rect 515 21 517 23
rect 511 20 517 21
rect 574 31 578 35
rect 613 39 617 45
rect 613 35 624 39
rect 574 27 598 31
rect 594 24 598 27
rect 620 29 624 35
rect 620 27 621 29
rect 623 27 624 29
rect 620 25 624 27
rect 594 22 595 24
rect 597 22 598 24
rect 594 20 598 22
rect 605 21 611 22
rect 605 19 607 21
rect 609 19 611 21
rect 534 16 540 17
rect 534 14 536 16
rect 538 14 540 16
rect 534 13 540 14
rect 553 16 559 17
rect 553 14 555 16
rect 557 14 559 16
rect 553 13 559 14
rect 605 13 611 19
<< via1 >>
rect 89 51 91 53
rect 40 36 42 38
rect 98 51 100 53
rect 81 27 83 29
rect 106 27 108 29
rect 153 28 155 30
rect 203 51 205 53
rect 171 36 173 38
rect 212 51 214 53
rect 195 27 197 29
rect 267 43 269 45
rect 220 27 222 29
rect 333 52 335 54
rect 314 28 316 30
rect 331 28 333 30
rect 356 44 358 46
rect 380 36 382 38
rect 407 36 409 38
rect 438 28 440 30
rect 505 52 507 54
rect 481 43 483 45
rect 458 28 460 30
rect 506 28 508 30
rect 524 44 526 46
rect 566 28 568 30
<< labels >>
rlabel alu1 126 9 126 9 6 vss
rlabel alu1 126 73 126 73 6 vdd
rlabel alu1 74 73 74 73 6 vdd
rlabel alu1 74 9 74 9 6 vss
rlabel alu1 240 9 240 9 6 vss
rlabel alu1 240 73 240 73 6 vdd
rlabel alu1 268 33 268 33 1 sum
rlabel alu1 188 73 188 73 6 vdd
rlabel alu1 188 9 188 9 6 vss
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 74 36 74 36 1 a
rlabel via1 89 51 89 51 1 b
rlabel via1 205 52 205 52 1 cin
rlabel alu1 9 39 9 39 1 cout
rlabel alu1 299 9 299 9 4 vss
rlabel alu1 299 37 299 37 4 a
rlabel alu1 291 33 291 33 4 a
rlabel alu1 291 45 291 45 4 b
rlabel alu1 299 73 299 73 4 vdd
rlabel alu1 283 53 283 53 4 b
rlabel alu1 400 61 400 61 6 z
rlabel alu1 420 9 420 9 6 vss
rlabel alu1 420 73 420 73 6 vdd
rlabel via1 357 45 357 45 4 a0
rlabel alu1 365 41 365 41 4 a0
rlabel alu1 353 9 353 9 4 vss
rlabel alu1 341 37 341 37 4 a1
rlabel alu1 353 73 353 73 4 vdd
rlabel alu1 333 29 333 29 4 a1
rlabel alu1 487 9 487 9 6 vss
rlabel alu1 487 73 487 73 6 vdd
rlabel alu1 479 44 479 44 1 a2
rlabel alu1 475 39 475 39 1 a2
rlabel alu1 498 37 498 37 1 a3
rlabel alu1 503 28 503 28 1 a3
rlabel via1 507 53 507 53 1 s1
rlabel alu1 515 61 515 61 1 s1
rlabel via1 333 53 333 53 1 s1
rlabel alu1 325 61 325 61 1 s1
rlabel alu1 448 61 448 61 1 s0
rlabel alu1 541 9 541 9 6 vss
rlabel alu1 541 73 541 73 6 vdd
rlabel alu1 557 53 557 53 6 b
rlabel alu1 557 29 557 29 6 a
rlabel alu1 541 45 541 45 6 b
rlabel alu1 549 45 549 45 6 b
rlabel alu1 549 37 549 37 6 a
rlabel alu1 541 37 541 37 6 a
rlabel alu1 615 29 615 29 4 a
rlabel alu1 623 53 623 53 4 b
rlabel alu1 615 61 615 61 4 b
rlabel alu1 607 33 607 33 4 a
rlabel alu1 595 9 595 9 4 vss
rlabel alu1 595 73 595 73 4 vdd
<< end >>
