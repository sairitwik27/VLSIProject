magic
tech scmos
timestamp 1608808693
<< ab >>
rect -34 5 6 77
rect 7 5 149 77
rect 151 5 190 77
rect 194 5 234 77
rect 236 5 339 77
<< nwell >>
rect -39 37 341 82
<< pwell >>
rect -39 0 341 37
<< poly >>
rect -25 62 -23 66
rect -15 64 -13 69
rect -5 64 -3 69
rect 15 64 17 69
rect 25 64 27 69
rect 95 71 97 75
rect 35 62 37 66
rect 55 64 57 69
rect 65 64 67 69
rect -25 40 -23 44
rect -15 40 -13 51
rect -5 48 -3 51
rect 15 48 17 51
rect -5 46 1 48
rect -5 44 -3 46
rect -1 44 1 46
rect -5 42 1 44
rect 11 46 17 48
rect 11 44 13 46
rect 15 44 17 46
rect 11 42 17 44
rect -25 38 -19 40
rect -25 36 -23 38
rect -21 36 -19 38
rect -25 34 -19 36
rect -15 38 -9 40
rect -15 36 -13 38
rect -11 36 -9 38
rect -15 34 -9 36
rect -25 29 -23 34
rect -12 29 -10 34
rect -5 29 -3 42
rect 15 29 17 42
rect 25 40 27 51
rect 75 62 77 66
rect 55 48 57 51
rect 51 46 57 48
rect 51 44 53 46
rect 55 44 57 46
rect 35 40 37 44
rect 51 42 57 44
rect 21 38 27 40
rect 21 36 23 38
rect 25 36 27 38
rect 21 34 27 36
rect 31 38 37 40
rect 31 36 33 38
rect 35 36 37 38
rect 31 34 37 36
rect 22 29 24 34
rect 35 29 37 34
rect 55 29 57 42
rect 65 40 67 51
rect 131 71 133 75
rect 105 62 107 66
rect 115 62 117 66
rect 160 64 162 69
rect 170 64 172 69
rect 252 71 254 75
rect 180 62 182 66
rect 203 62 205 66
rect 213 64 215 69
rect 223 64 225 69
rect 160 48 162 51
rect 142 46 148 48
rect 142 44 144 46
rect 146 44 148 46
rect 75 40 77 44
rect 61 38 67 40
rect 61 36 63 38
rect 65 36 67 38
rect 61 34 67 36
rect 71 38 77 40
rect 71 36 73 38
rect 75 36 77 38
rect 71 34 77 36
rect 95 41 97 44
rect 95 39 101 41
rect 95 37 97 39
rect 99 37 101 39
rect 95 35 101 37
rect 105 40 107 44
rect 115 41 117 44
rect 131 41 133 44
rect 142 42 148 44
rect 156 46 162 48
rect 156 44 158 46
rect 160 44 162 46
rect 156 42 162 44
rect 142 41 144 42
rect 105 38 111 40
rect 115 39 125 41
rect 131 39 144 41
rect 105 36 107 38
rect 109 36 111 38
rect 62 29 64 34
rect 75 29 77 34
rect -25 16 -23 20
rect -12 13 -10 18
rect -5 13 -3 18
rect 15 13 17 18
rect 22 13 24 18
rect 35 16 37 20
rect 96 26 98 35
rect 105 34 111 36
rect 123 35 125 39
rect 105 31 107 34
rect 103 29 107 31
rect 123 33 132 35
rect 123 31 128 33
rect 130 31 132 33
rect 139 31 141 39
rect 103 26 105 29
rect 113 26 115 30
rect 123 29 132 31
rect 123 26 125 29
rect 55 13 57 18
rect 62 13 64 18
rect 75 16 77 20
rect 160 29 162 42
rect 170 40 172 51
rect 180 40 182 44
rect 166 38 172 40
rect 166 36 168 38
rect 170 36 172 38
rect 166 34 172 36
rect 176 38 182 40
rect 176 36 178 38
rect 180 36 182 38
rect 176 34 182 36
rect 167 29 169 34
rect 180 29 182 34
rect 203 40 205 44
rect 213 40 215 51
rect 223 48 225 51
rect 223 46 229 48
rect 223 44 225 46
rect 227 44 229 46
rect 223 42 229 44
rect 237 46 243 48
rect 237 44 239 46
rect 241 44 243 46
rect 288 71 290 75
rect 268 62 270 66
rect 278 62 280 66
rect 308 62 310 66
rect 318 64 320 69
rect 328 64 330 69
rect 237 42 243 44
rect 203 38 209 40
rect 203 36 205 38
rect 207 36 209 38
rect 203 34 209 36
rect 213 38 219 40
rect 213 36 215 38
rect 217 36 219 38
rect 213 34 219 36
rect 203 29 205 34
rect 216 29 218 34
rect 223 29 225 42
rect 241 41 243 42
rect 252 41 254 44
rect 268 41 270 44
rect 241 39 254 41
rect 260 39 270 41
rect 278 40 280 44
rect 288 41 290 44
rect 244 31 246 39
rect 260 35 262 39
rect 253 33 262 35
rect 274 38 280 40
rect 274 36 276 38
rect 278 36 280 38
rect 274 34 280 36
rect 284 39 290 41
rect 284 37 286 39
rect 288 37 290 39
rect 284 35 290 37
rect 308 40 310 44
rect 318 40 320 51
rect 328 48 330 51
rect 328 46 334 48
rect 328 44 330 46
rect 332 44 334 46
rect 328 42 334 44
rect 308 38 314 40
rect 308 36 310 38
rect 312 36 314 38
rect 253 31 255 33
rect 257 31 262 33
rect 139 19 141 22
rect 136 17 141 19
rect 96 9 98 14
rect 103 9 105 14
rect 113 9 115 17
rect 123 13 125 17
rect 136 9 138 17
rect 113 7 138 9
rect 160 13 162 18
rect 167 13 169 18
rect 180 16 182 20
rect 203 16 205 20
rect 253 29 262 31
rect 278 31 280 34
rect 260 26 262 29
rect 270 26 272 30
rect 278 29 282 31
rect 280 26 282 29
rect 287 26 289 35
rect 308 34 314 36
rect 318 38 324 40
rect 318 36 320 38
rect 322 36 324 38
rect 318 34 324 36
rect 308 29 310 34
rect 321 29 323 34
rect 328 29 330 42
rect 244 19 246 22
rect 216 13 218 18
rect 223 13 225 18
rect 244 17 249 19
rect 247 9 249 17
rect 260 13 262 17
rect 270 9 272 17
rect 308 16 310 20
rect 280 9 282 14
rect 287 9 289 14
rect 247 7 272 9
rect 321 13 323 18
rect 328 13 330 18
<< ndif >>
rect -30 26 -25 29
rect -32 24 -25 26
rect -32 22 -30 24
rect -28 22 -25 24
rect -32 20 -25 22
rect -23 20 -12 29
rect -21 18 -12 20
rect -10 18 -5 29
rect -3 24 2 29
rect 10 24 15 29
rect -3 22 4 24
rect -3 20 0 22
rect 2 20 4 22
rect -3 18 4 20
rect 8 22 15 24
rect 8 20 10 22
rect 12 20 15 22
rect 8 18 15 20
rect 17 18 22 29
rect 24 20 35 29
rect 37 26 42 29
rect 37 24 44 26
rect 50 24 55 29
rect 37 22 40 24
rect 42 22 44 24
rect 37 20 44 22
rect 48 22 55 24
rect 48 20 50 22
rect 52 20 55 22
rect 24 18 33 20
rect -21 12 -14 18
rect -21 10 -19 12
rect -17 10 -14 12
rect -21 8 -14 10
rect 26 12 33 18
rect 48 18 55 20
rect 57 18 62 29
rect 64 20 75 29
rect 77 26 82 29
rect 134 26 139 31
rect 77 24 84 26
rect 77 22 80 24
rect 82 22 84 24
rect 77 20 84 22
rect 64 18 73 20
rect 26 10 29 12
rect 31 10 33 12
rect 26 8 33 10
rect 66 12 73 18
rect 88 14 96 26
rect 98 14 103 26
rect 105 22 113 26
rect 105 20 108 22
rect 110 20 113 22
rect 105 17 113 20
rect 115 24 123 26
rect 115 22 118 24
rect 120 22 123 24
rect 115 17 123 22
rect 125 22 139 26
rect 141 29 148 31
rect 237 29 244 31
rect 141 27 144 29
rect 146 27 148 29
rect 141 25 148 27
rect 141 22 146 25
rect 155 24 160 29
rect 153 22 160 24
rect 125 21 134 22
rect 125 19 130 21
rect 132 19 134 21
rect 125 17 134 19
rect 153 20 155 22
rect 157 20 160 22
rect 153 18 160 20
rect 162 18 167 29
rect 169 20 180 29
rect 182 26 187 29
rect 198 26 203 29
rect 182 24 189 26
rect 182 22 185 24
rect 187 22 189 24
rect 182 20 189 22
rect 196 24 203 26
rect 196 22 198 24
rect 200 22 203 24
rect 196 20 203 22
rect 205 20 216 29
rect 169 18 178 20
rect 105 14 110 17
rect 66 10 69 12
rect 71 10 73 12
rect 66 8 73 10
rect 88 12 94 14
rect 88 10 90 12
rect 92 10 94 12
rect 88 8 94 10
rect 171 12 178 18
rect 207 18 216 20
rect 218 18 223 29
rect 225 24 230 29
rect 237 27 239 29
rect 241 27 244 29
rect 237 25 244 27
rect 225 22 232 24
rect 239 22 244 25
rect 246 26 251 31
rect 303 26 308 29
rect 246 22 260 26
rect 225 20 228 22
rect 230 20 232 22
rect 225 18 232 20
rect 251 21 260 22
rect 251 19 253 21
rect 255 19 260 21
rect 171 10 174 12
rect 176 10 178 12
rect 171 8 178 10
rect 207 12 214 18
rect 251 17 260 19
rect 262 24 270 26
rect 262 22 265 24
rect 267 22 270 24
rect 262 17 270 22
rect 272 22 280 26
rect 272 20 275 22
rect 277 20 280 22
rect 272 17 280 20
rect 207 10 209 12
rect 211 10 214 12
rect 207 8 214 10
rect 275 14 280 17
rect 282 14 287 26
rect 289 14 297 26
rect 301 24 308 26
rect 301 22 303 24
rect 305 22 308 24
rect 301 20 308 22
rect 310 20 321 29
rect 312 18 321 20
rect 323 18 328 29
rect 330 24 335 29
rect 330 22 337 24
rect 330 20 333 22
rect 335 20 337 22
rect 330 18 337 20
rect 291 12 297 14
rect 291 10 293 12
rect 295 10 297 12
rect 291 8 297 10
rect 312 12 319 18
rect 312 10 314 12
rect 316 10 319 12
rect 312 8 319 10
<< pdif >>
rect -21 62 -15 64
rect -30 57 -25 62
rect -32 55 -25 57
rect -32 53 -30 55
rect -28 53 -25 55
rect -32 48 -25 53
rect -32 46 -30 48
rect -28 46 -25 48
rect -32 44 -25 46
rect -23 60 -15 62
rect -23 58 -20 60
rect -18 58 -15 60
rect -23 51 -15 58
rect -13 62 -5 64
rect -13 60 -10 62
rect -8 60 -5 62
rect -13 55 -5 60
rect -13 53 -10 55
rect -8 53 -5 55
rect -13 51 -5 53
rect -3 62 4 64
rect -3 60 0 62
rect 2 60 4 62
rect -3 51 4 60
rect 8 62 15 64
rect 8 60 10 62
rect 12 60 15 62
rect 8 51 15 60
rect 17 62 25 64
rect 17 60 20 62
rect 22 60 25 62
rect 17 55 25 60
rect 17 53 20 55
rect 22 53 25 55
rect 17 51 25 53
rect 27 62 33 64
rect 48 62 55 64
rect 27 60 35 62
rect 27 58 30 60
rect 32 58 35 60
rect 27 51 35 58
rect -23 44 -17 51
rect 29 44 35 51
rect 37 57 42 62
rect 48 60 50 62
rect 52 60 55 62
rect 37 55 44 57
rect 37 53 40 55
rect 42 53 44 55
rect 37 48 44 53
rect 48 51 55 60
rect 57 62 65 64
rect 57 60 60 62
rect 62 60 65 62
rect 57 55 65 60
rect 57 53 60 55
rect 62 53 65 55
rect 57 51 65 53
rect 67 62 73 64
rect 90 65 95 71
rect 88 63 95 65
rect 67 60 75 62
rect 67 58 70 60
rect 72 58 75 60
rect 67 51 75 58
rect 37 46 40 48
rect 42 46 44 48
rect 37 44 44 46
rect 69 44 75 51
rect 77 57 82 62
rect 88 61 90 63
rect 92 61 95 63
rect 88 59 95 61
rect 77 55 84 57
rect 77 53 80 55
rect 82 53 84 55
rect 77 48 84 53
rect 77 46 80 48
rect 82 46 84 48
rect 77 44 84 46
rect 90 44 95 59
rect 97 62 102 71
rect 119 69 131 71
rect 119 67 126 69
rect 128 67 131 69
rect 119 62 131 67
rect 97 55 105 62
rect 97 53 100 55
rect 102 53 105 55
rect 97 44 105 53
rect 107 55 115 62
rect 107 53 110 55
rect 112 53 115 55
rect 107 48 115 53
rect 107 46 110 48
rect 112 46 115 48
rect 107 44 115 46
rect 117 60 126 62
rect 128 60 131 62
rect 117 44 131 60
rect 133 50 138 71
rect 153 62 160 64
rect 153 60 155 62
rect 157 60 160 62
rect 153 51 160 60
rect 162 62 170 64
rect 162 60 165 62
rect 167 60 170 62
rect 162 55 170 60
rect 162 53 165 55
rect 167 53 170 55
rect 162 51 170 53
rect 172 62 178 64
rect 207 62 213 64
rect 172 60 180 62
rect 172 58 175 60
rect 177 58 180 60
rect 172 51 180 58
rect 133 48 140 50
rect 133 46 136 48
rect 138 46 140 48
rect 133 44 140 46
rect 174 44 180 51
rect 182 57 187 62
rect 198 57 203 62
rect 182 55 189 57
rect 182 53 185 55
rect 187 53 189 55
rect 182 48 189 53
rect 182 46 185 48
rect 187 46 189 48
rect 182 44 189 46
rect 196 55 203 57
rect 196 53 198 55
rect 200 53 203 55
rect 196 48 203 53
rect 196 46 198 48
rect 200 46 203 48
rect 196 44 203 46
rect 205 60 213 62
rect 205 58 208 60
rect 210 58 213 60
rect 205 51 213 58
rect 215 62 223 64
rect 215 60 218 62
rect 220 60 223 62
rect 215 55 223 60
rect 215 53 218 55
rect 220 53 223 55
rect 215 51 223 53
rect 225 62 232 64
rect 225 60 228 62
rect 230 60 232 62
rect 225 51 232 60
rect 205 44 211 51
rect 247 50 252 71
rect 245 48 252 50
rect 245 46 247 48
rect 249 46 252 48
rect 245 44 252 46
rect 254 69 266 71
rect 254 67 257 69
rect 259 67 266 69
rect 254 62 266 67
rect 283 62 288 71
rect 254 60 257 62
rect 259 60 268 62
rect 254 44 268 60
rect 270 55 278 62
rect 270 53 273 55
rect 275 53 278 55
rect 270 48 278 53
rect 270 46 273 48
rect 275 46 278 48
rect 270 44 278 46
rect 280 55 288 62
rect 280 53 283 55
rect 285 53 288 55
rect 280 44 288 53
rect 290 65 295 71
rect 290 63 297 65
rect 290 61 293 63
rect 295 61 297 63
rect 312 62 318 64
rect 290 59 297 61
rect 290 44 295 59
rect 303 57 308 62
rect 301 55 308 57
rect 301 53 303 55
rect 305 53 308 55
rect 301 48 308 53
rect 301 46 303 48
rect 305 46 308 48
rect 301 44 308 46
rect 310 60 318 62
rect 310 58 313 60
rect 315 58 318 60
rect 310 51 318 58
rect 320 62 328 64
rect 320 60 323 62
rect 325 60 328 62
rect 320 55 328 60
rect 320 53 323 55
rect 325 53 328 55
rect 320 51 328 53
rect 330 62 337 64
rect 330 60 333 62
rect 335 60 337 62
rect 330 51 337 60
rect 310 44 316 51
<< alu1 >>
rect -36 72 341 77
rect -36 70 -29 72
rect -27 70 39 72
rect 41 70 79 72
rect 81 70 110 72
rect 112 70 184 72
rect 186 70 199 72
rect 201 70 273 72
rect 275 70 304 72
rect 306 70 341 72
rect -36 69 341 70
rect -32 55 -27 57
rect -32 53 -30 55
rect -28 53 -27 55
rect -32 48 -27 53
rect -32 46 -30 48
rect -28 46 -27 48
rect -32 44 -27 46
rect -32 24 -28 44
rect 0 47 4 56
rect -9 46 4 47
rect -9 44 -3 46
rect -1 44 4 46
rect -9 43 4 44
rect 8 47 12 56
rect 39 55 44 57
rect 8 46 21 47
rect 8 44 13 46
rect 15 44 21 46
rect 8 43 21 44
rect -17 38 -3 39
rect -17 36 -13 38
rect -11 36 -3 38
rect -17 35 -3 36
rect -32 22 -30 24
rect -28 22 -20 24
rect -32 18 -20 22
rect -8 26 -3 35
rect 15 38 29 39
rect 15 36 23 38
rect 25 36 29 38
rect 15 35 29 36
rect 39 53 40 55
rect 42 53 44 55
rect 39 52 44 53
rect 39 50 40 52
rect 42 50 44 52
rect 39 48 44 50
rect 39 46 40 48
rect 42 46 44 48
rect 39 44 44 46
rect 15 26 20 35
rect 40 24 44 44
rect 48 47 52 56
rect 79 55 84 57
rect 48 46 61 47
rect 48 44 53 46
rect 55 44 61 46
rect 48 43 61 44
rect 55 38 69 39
rect 55 36 63 38
rect 65 36 69 38
rect 55 35 69 36
rect 79 53 80 55
rect 82 53 84 55
rect 79 48 84 53
rect 79 46 80 48
rect 82 46 84 48
rect 79 44 84 46
rect 55 26 60 35
rect 80 29 84 44
rect 80 27 81 29
rect 83 27 84 29
rect 32 22 40 24
rect 42 22 44 24
rect 80 24 84 27
rect 32 18 44 22
rect 72 22 80 24
rect 82 22 84 24
rect 72 18 84 22
rect 88 55 104 56
rect 88 53 100 55
rect 102 53 104 55
rect 88 51 104 53
rect 88 23 92 51
rect 136 58 148 64
rect 143 52 148 58
rect 143 50 144 52
rect 146 50 148 52
rect 143 49 148 50
rect 153 49 157 56
rect 184 55 189 57
rect 127 33 132 40
rect 143 47 157 49
rect 143 46 166 47
rect 143 44 144 46
rect 146 44 158 46
rect 160 44 166 46
rect 143 43 149 44
rect 153 43 166 44
rect 143 42 148 43
rect 127 31 128 33
rect 130 32 132 33
rect 130 31 140 32
rect 127 29 140 31
rect 127 27 135 29
rect 137 27 140 29
rect 127 26 140 27
rect 160 38 174 39
rect 160 36 168 38
rect 170 36 174 38
rect 160 35 174 36
rect 184 53 185 55
rect 187 53 189 55
rect 184 48 189 53
rect 184 46 185 48
rect 187 46 189 48
rect 184 45 189 46
rect 184 44 186 45
rect 160 29 165 35
rect 160 27 162 29
rect 164 27 165 29
rect 160 26 165 27
rect 185 43 186 44
rect 188 43 189 45
rect 88 22 112 23
rect 88 20 108 22
rect 110 20 112 22
rect 185 24 189 43
rect 88 19 112 20
rect 177 22 185 24
rect 187 22 189 24
rect 177 18 189 22
rect 196 55 201 57
rect 196 53 198 55
rect 200 53 201 55
rect 237 58 249 64
rect 196 48 201 53
rect 196 46 198 48
rect 200 46 201 48
rect 196 44 201 46
rect 196 24 200 44
rect 228 49 232 56
rect 237 49 242 58
rect 228 47 242 49
rect 219 46 242 47
rect 219 44 220 46
rect 222 44 225 46
rect 227 44 239 46
rect 241 44 242 46
rect 219 43 232 44
rect 236 43 242 44
rect 237 42 242 43
rect 211 38 225 39
rect 211 36 215 38
rect 217 36 225 38
rect 211 35 225 36
rect 196 22 198 24
rect 200 22 208 24
rect 196 18 208 22
rect 220 29 225 35
rect 220 27 221 29
rect 223 27 225 29
rect 220 26 225 27
rect 253 33 258 40
rect 281 55 297 56
rect 281 53 283 55
rect 285 53 297 55
rect 281 51 297 53
rect 253 32 255 33
rect 245 31 255 32
rect 257 31 258 33
rect 245 29 258 31
rect 245 27 248 29
rect 250 27 258 29
rect 245 26 258 27
rect 293 23 297 51
rect 273 22 297 23
rect 273 20 275 22
rect 277 20 297 22
rect 273 19 297 20
rect 301 55 306 57
rect 301 53 303 55
rect 305 53 306 55
rect 301 48 306 53
rect 301 46 303 48
rect 305 46 306 48
rect 301 44 306 46
rect 301 29 305 44
rect 301 27 302 29
rect 304 27 305 29
rect 333 47 337 56
rect 324 46 337 47
rect 324 44 330 46
rect 332 44 337 46
rect 324 43 337 44
rect 316 38 330 39
rect 316 36 320 38
rect 322 36 330 38
rect 316 35 330 36
rect 301 24 305 27
rect 301 22 303 24
rect 305 22 313 24
rect 301 18 313 22
rect 325 26 330 35
rect -36 12 341 13
rect -36 10 -29 12
rect -27 10 -19 12
rect -17 10 29 12
rect 31 10 39 12
rect 41 10 69 12
rect 71 10 79 12
rect 81 10 90 12
rect 92 10 143 12
rect 145 10 174 12
rect 176 10 184 12
rect 186 10 199 12
rect 201 10 209 12
rect 211 10 240 12
rect 242 10 293 12
rect 295 10 304 12
rect 306 10 314 12
rect 316 10 341 12
rect -36 5 341 10
<< alu2 >>
rect 39 52 148 54
rect 39 50 40 52
rect 42 50 144 52
rect 146 50 148 52
rect 39 49 148 50
rect 185 46 231 47
rect 185 45 220 46
rect 185 43 186 45
rect 188 44 220 45
rect 222 44 231 46
rect 188 43 231 44
rect 185 42 189 43
rect 80 29 165 30
rect 80 27 81 29
rect 83 27 135 29
rect 137 27 162 29
rect 164 27 165 29
rect 80 26 165 27
rect 220 29 305 30
rect 220 27 221 29
rect 223 27 248 29
rect 250 27 302 29
rect 304 27 305 29
rect 220 26 305 27
<< ptie >>
rect -31 12 -25 14
rect -31 10 -29 12
rect -27 10 -25 12
rect -31 8 -25 10
rect 37 12 43 14
rect 37 10 39 12
rect 41 10 43 12
rect 37 8 43 10
rect 77 12 83 14
rect 77 10 79 12
rect 81 10 83 12
rect 77 8 83 10
rect 141 12 147 14
rect 141 10 143 12
rect 145 10 147 12
rect 141 8 147 10
rect 182 12 188 14
rect 182 10 184 12
rect 186 10 188 12
rect 182 8 188 10
rect 197 12 203 14
rect 197 10 199 12
rect 201 10 203 12
rect 197 8 203 10
rect 238 12 244 14
rect 238 10 240 12
rect 242 10 244 12
rect 238 8 244 10
rect 302 12 308 14
rect 302 10 304 12
rect 306 10 308 12
rect 302 8 308 10
<< ntie >>
rect -31 72 -25 74
rect -31 70 -29 72
rect -27 70 -25 72
rect -31 68 -25 70
rect 37 72 43 74
rect 37 70 39 72
rect 41 70 43 72
rect 37 68 43 70
rect 77 72 83 74
rect 77 70 79 72
rect 81 70 83 72
rect 108 72 114 74
rect 77 68 83 70
rect 108 70 110 72
rect 112 70 114 72
rect 182 72 188 74
rect 108 68 114 70
rect 182 70 184 72
rect 186 70 188 72
rect 182 68 188 70
rect 197 72 203 74
rect 197 70 199 72
rect 201 70 203 72
rect 271 72 277 74
rect 197 68 203 70
rect 271 70 273 72
rect 275 70 277 72
rect 302 72 308 74
rect 271 68 277 70
rect 302 70 304 72
rect 306 70 308 72
rect 302 68 308 70
<< nmos >>
rect -25 20 -23 29
rect -12 18 -10 29
rect -5 18 -3 29
rect 15 18 17 29
rect 22 18 24 29
rect 35 20 37 29
rect 55 18 57 29
rect 62 18 64 29
rect 75 20 77 29
rect 96 14 98 26
rect 103 14 105 26
rect 113 17 115 26
rect 123 17 125 26
rect 139 22 141 31
rect 160 18 162 29
rect 167 18 169 29
rect 180 20 182 29
rect 203 20 205 29
rect 216 18 218 29
rect 223 18 225 29
rect 244 22 246 31
rect 260 17 262 26
rect 270 17 272 26
rect 280 14 282 26
rect 287 14 289 26
rect 308 20 310 29
rect 321 18 323 29
rect 328 18 330 29
<< pmos >>
rect -25 44 -23 62
rect -15 51 -13 64
rect -5 51 -3 64
rect 15 51 17 64
rect 25 51 27 64
rect 35 44 37 62
rect 55 51 57 64
rect 65 51 67 64
rect 75 44 77 62
rect 95 44 97 71
rect 105 44 107 62
rect 115 44 117 62
rect 131 44 133 71
rect 160 51 162 64
rect 170 51 172 64
rect 180 44 182 62
rect 203 44 205 62
rect 213 51 215 64
rect 223 51 225 64
rect 252 44 254 71
rect 268 44 270 62
rect 278 44 280 62
rect 288 44 290 71
rect 308 44 310 62
rect 318 51 320 64
rect 328 51 330 64
<< polyct0 >>
rect -23 36 -21 38
rect 33 36 35 38
rect 73 36 75 38
rect 97 37 99 39
rect 107 36 109 38
rect 178 36 180 38
rect 205 36 207 38
rect 276 36 278 38
rect 286 37 288 39
rect 310 36 312 38
<< polyct1 >>
rect -3 44 -1 46
rect 13 44 15 46
rect -13 36 -11 38
rect 53 44 55 46
rect 23 36 25 38
rect 144 44 146 46
rect 63 36 65 38
rect 158 44 160 46
rect 128 31 130 33
rect 168 36 170 38
rect 225 44 227 46
rect 239 44 241 46
rect 215 36 217 38
rect 330 44 332 46
rect 255 31 257 33
rect 320 36 322 38
<< ndifct0 >>
rect 0 20 2 22
rect 10 20 12 22
rect 50 20 52 22
rect 118 22 120 24
rect 144 27 146 29
rect 130 19 132 21
rect 155 20 157 22
rect 239 27 241 29
rect 228 20 230 22
rect 253 19 255 21
rect 265 22 267 24
rect 333 20 335 22
<< ndifct1 >>
rect -30 22 -28 24
rect 40 22 42 24
rect -19 10 -17 12
rect 80 22 82 24
rect 29 10 31 12
rect 108 20 110 22
rect 185 22 187 24
rect 198 22 200 24
rect 69 10 71 12
rect 90 10 92 12
rect 174 10 176 12
rect 275 20 277 22
rect 209 10 211 12
rect 303 22 305 24
rect 293 10 295 12
rect 314 10 316 12
<< ntiect1 >>
rect -29 70 -27 72
rect 39 70 41 72
rect 79 70 81 72
rect 110 70 112 72
rect 184 70 186 72
rect 199 70 201 72
rect 273 70 275 72
rect 304 70 306 72
<< ptiect1 >>
rect -29 10 -27 12
rect 39 10 41 12
rect 79 10 81 12
rect 143 10 145 12
rect 184 10 186 12
rect 199 10 201 12
rect 240 10 242 12
rect 304 10 306 12
<< pdifct0 >>
rect -20 58 -18 60
rect -10 60 -8 62
rect -10 53 -8 55
rect 0 60 2 62
rect 10 60 12 62
rect 20 60 22 62
rect 20 53 22 55
rect 30 58 32 60
rect 50 60 52 62
rect 60 60 62 62
rect 60 53 62 55
rect 70 58 72 60
rect 90 61 92 63
rect 126 67 128 69
rect 110 53 112 55
rect 110 46 112 48
rect 126 60 128 62
rect 155 60 157 62
rect 165 60 167 62
rect 165 53 167 55
rect 175 58 177 60
rect 136 46 138 48
rect 208 58 210 60
rect 218 60 220 62
rect 218 53 220 55
rect 228 60 230 62
rect 247 46 249 48
rect 257 67 259 69
rect 257 60 259 62
rect 273 53 275 55
rect 273 46 275 48
rect 293 61 295 63
rect 313 58 315 60
rect 323 60 325 62
rect 323 53 325 55
rect 333 60 335 62
<< pdifct1 >>
rect -30 53 -28 55
rect -30 46 -28 48
rect 40 53 42 55
rect 40 46 42 48
rect 80 53 82 55
rect 80 46 82 48
rect 100 53 102 55
rect 185 53 187 55
rect 185 46 187 48
rect 198 53 200 55
rect 198 46 200 48
rect 283 53 285 55
rect 303 53 305 55
rect 303 46 305 48
<< alu0 >>
rect -22 60 -16 69
rect -22 58 -20 60
rect -18 58 -16 60
rect -22 57 -16 58
rect -11 62 -7 64
rect -11 60 -10 62
rect -8 60 -7 62
rect -11 55 -7 60
rect -2 62 4 69
rect -2 60 0 62
rect 2 60 4 62
rect -2 59 4 60
rect 8 62 14 69
rect 8 60 10 62
rect 12 60 14 62
rect 8 59 14 60
rect 19 62 23 64
rect 19 60 20 62
rect 22 60 23 62
rect -11 54 -10 55
rect -24 53 -10 54
rect -8 53 -7 55
rect -24 50 -7 53
rect -24 38 -20 50
rect 19 55 23 60
rect 28 60 34 69
rect 28 58 30 60
rect 32 58 34 60
rect 48 62 54 69
rect 48 60 50 62
rect 52 60 54 62
rect 48 59 54 60
rect 59 62 63 64
rect 59 60 60 62
rect 62 60 63 62
rect 28 57 34 58
rect 19 53 20 55
rect 22 54 23 55
rect 22 53 36 54
rect 19 50 36 53
rect -24 36 -23 38
rect -21 36 -20 38
rect -24 31 -20 36
rect -24 27 -12 31
rect -28 24 -27 26
rect -16 23 -12 27
rect 32 38 36 50
rect 32 36 33 38
rect 35 36 36 38
rect 32 31 36 36
rect 24 27 36 31
rect 24 23 28 27
rect 39 24 40 26
rect 59 55 63 60
rect 68 60 74 69
rect 125 67 126 69
rect 128 67 129 69
rect 88 63 121 64
rect 88 61 90 63
rect 92 61 121 63
rect 88 60 121 61
rect 68 58 70 60
rect 72 58 74 60
rect 68 57 74 58
rect 59 53 60 55
rect 62 54 63 55
rect 62 53 76 54
rect 59 50 76 53
rect 72 38 76 50
rect 72 36 73 38
rect 75 36 76 38
rect 72 31 76 36
rect 64 27 76 31
rect -16 22 4 23
rect -16 20 0 22
rect 2 20 4 22
rect -16 19 4 20
rect 8 22 28 23
rect 8 20 10 22
rect 12 20 28 22
rect 8 19 28 20
rect 64 23 68 27
rect 79 24 80 26
rect 48 22 68 23
rect 48 20 50 22
rect 52 20 68 22
rect 48 19 68 20
rect 109 55 113 57
rect 109 53 110 55
rect 112 53 113 55
rect 109 48 113 53
rect 109 47 110 48
rect 97 46 110 47
rect 112 46 113 48
rect 97 43 113 46
rect 117 49 121 60
rect 125 62 129 67
rect 125 60 126 62
rect 128 60 129 62
rect 125 58 129 60
rect 153 62 159 69
rect 153 60 155 62
rect 157 60 159 62
rect 153 59 159 60
rect 164 62 168 64
rect 164 60 165 62
rect 167 60 168 62
rect 164 55 168 60
rect 173 60 179 69
rect 173 58 175 60
rect 177 58 179 60
rect 173 57 179 58
rect 206 60 212 69
rect 206 58 208 60
rect 210 58 212 60
rect 206 57 212 58
rect 217 62 221 64
rect 217 60 218 62
rect 220 60 221 62
rect 164 53 165 55
rect 167 54 168 55
rect 167 53 181 54
rect 164 50 181 53
rect 117 48 140 49
rect 117 46 136 48
rect 138 46 140 48
rect 117 45 140 46
rect 97 41 101 43
rect 96 39 101 41
rect 117 39 121 45
rect 96 37 97 39
rect 99 37 101 39
rect 96 35 101 37
rect 105 38 121 39
rect 105 36 107 38
rect 109 36 121 38
rect 105 35 121 36
rect 97 31 101 35
rect 136 39 140 45
rect 136 35 147 39
rect 97 27 121 31
rect 117 24 121 27
rect 143 29 147 35
rect 143 27 144 29
rect 146 27 147 29
rect 143 25 147 27
rect 177 38 181 50
rect 177 36 178 38
rect 180 36 181 38
rect 177 31 181 36
rect 169 27 181 31
rect 117 22 118 24
rect 120 22 121 24
rect 169 23 173 27
rect 184 24 185 26
rect 153 22 173 23
rect 117 20 121 22
rect 128 21 134 22
rect 128 19 130 21
rect 132 19 134 21
rect 153 20 155 22
rect 157 20 173 22
rect 153 19 173 20
rect 128 13 134 19
rect 217 55 221 60
rect 226 62 232 69
rect 256 67 257 69
rect 259 67 260 69
rect 226 60 228 62
rect 230 60 232 62
rect 226 59 232 60
rect 256 62 260 67
rect 256 60 257 62
rect 259 60 260 62
rect 256 58 260 60
rect 264 63 297 64
rect 264 61 293 63
rect 295 61 297 63
rect 264 60 297 61
rect 311 60 317 69
rect 217 54 218 55
rect 204 53 218 54
rect 220 53 221 55
rect 204 50 221 53
rect 204 38 208 50
rect 264 49 268 60
rect 311 58 313 60
rect 315 58 317 60
rect 311 57 317 58
rect 322 62 326 64
rect 322 60 323 62
rect 325 60 326 62
rect 245 48 268 49
rect 245 46 247 48
rect 249 46 268 48
rect 245 45 268 46
rect 245 39 249 45
rect 204 36 205 38
rect 207 36 208 38
rect 204 31 208 36
rect 204 27 216 31
rect 200 24 201 26
rect 212 23 216 27
rect 238 35 249 39
rect 238 29 242 35
rect 264 39 268 45
rect 272 55 276 57
rect 272 53 273 55
rect 275 53 276 55
rect 272 48 276 53
rect 272 46 273 48
rect 275 47 276 48
rect 275 46 288 47
rect 272 43 288 46
rect 284 41 288 43
rect 284 39 289 41
rect 264 38 280 39
rect 264 36 276 38
rect 278 36 280 38
rect 264 35 280 36
rect 284 37 286 39
rect 288 37 289 39
rect 284 35 289 37
rect 238 27 239 29
rect 241 27 242 29
rect 238 25 242 27
rect 284 31 288 35
rect 264 27 288 31
rect 264 24 268 27
rect 212 22 232 23
rect 264 22 265 24
rect 267 22 268 24
rect 212 20 228 22
rect 230 20 232 22
rect 212 19 232 20
rect 251 21 257 22
rect 251 19 253 21
rect 255 19 257 21
rect 264 20 268 22
rect 322 55 326 60
rect 331 62 337 69
rect 331 60 333 62
rect 335 60 337 62
rect 331 59 337 60
rect 322 54 323 55
rect 309 53 323 54
rect 325 53 326 55
rect 309 50 326 53
rect 309 38 313 50
rect 309 36 310 38
rect 312 36 313 38
rect 309 31 313 36
rect 309 27 321 31
rect 305 24 306 26
rect 251 13 257 19
rect 317 23 321 27
rect 317 22 337 23
rect 317 20 333 22
rect 335 20 337 22
rect 317 19 337 20
<< via1 >>
rect 40 50 42 52
rect 81 27 83 29
rect 144 50 146 52
rect 135 27 137 29
rect 162 27 164 29
rect 186 43 188 45
rect 220 44 222 46
rect 221 27 223 29
rect 248 27 250 29
rect 302 27 304 29
<< labels >>
rlabel alu1 238 73 238 73 1 Vdd
rlabel alu1 214 73 214 73 6 vdd
rlabel alu1 236 8 236 8 1 Vss
rlabel alu1 149 8 149 8 1 Vss
rlabel alu1 171 73 171 73 4 vdd
rlabel alu1 147 73 147 73 1 Vdd
rlabel alu1 66 9 66 9 4 vss
rlabel alu1 66 73 66 73 4 vdd
rlabel alu1 26 73 26 73 4 vdd
rlabel alu1 26 9 26 9 4 vss
rlabel alu1 319 73 319 73 6 vdd
rlabel alu1 319 9 319 9 6 vss
rlabel alu1 50 53 50 53 1 b0
rlabel alu1 58 33 58 33 1 a1
rlabel alu1 42 37 42 37 1 z1
rlabel alu1 18 33 18 33 1 a0
rlabel alu1 18 45 18 45 1 b1
rlabel alu1 90 40 90 40 1 p1
rlabel alu1 327 33 327 33 1 a1
rlabel alu1 335 53 335 53 1 b1
rlabel alu1 295 40 295 40 1 p2
rlabel alu1 198 35 198 35 1 p3
rlabel alu1 -14 73 -14 73 6 vdd
rlabel alu1 -14 9 -14 9 6 vss
rlabel alu1 2 53 2 53 1 b0
rlabel alu1 -6 33 -6 33 1 a0
rlabel alu1 -30 37 -30 37 1 p0
<< end >>
