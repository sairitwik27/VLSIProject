magic
tech scmos
timestamp 1608981221
<< ab >>
rect 4 410 52 418
rect 13 345 52 410
rect 54 345 90 418
rect 13 282 50 345
rect 4 274 50 282
rect 52 274 90 345
rect 92 410 97 418
rect 92 354 94 410
rect 92 345 97 354
rect 99 345 162 418
rect 164 386 202 418
rect 486 412 534 420
rect 164 345 211 386
rect 92 274 132 345
rect 134 274 197 345
rect 202 306 211 345
rect 495 347 534 412
rect 536 347 572 420
rect 495 284 532 347
rect 486 276 532 284
rect 534 276 572 347
rect 574 412 579 420
rect 574 356 576 412
rect 574 347 579 356
rect 581 347 644 420
rect 646 412 739 420
rect 646 388 684 412
rect 646 356 693 388
rect 700 356 739 412
rect 646 347 739 356
rect 741 347 777 420
rect 574 276 614 347
rect 616 276 679 347
rect 684 340 737 347
rect 684 308 693 340
rect 700 284 737 340
rect 681 276 737 284
rect 739 276 777 347
rect 779 412 784 420
rect 779 356 781 412
rect 779 347 784 356
rect 786 347 849 420
rect 851 388 889 420
rect 851 347 898 388
rect 779 276 819 347
rect 821 276 884 347
rect 889 308 898 347
rect 1012 294 1060 302
rect -1 158 79 230
rect 81 158 184 230
rect 186 158 329 230
rect 331 158 434 230
rect 436 158 579 230
rect 581 158 684 230
rect 686 158 829 230
rect 831 158 934 230
rect 936 158 999 230
rect 1021 229 1060 294
rect 1062 229 1098 302
rect 1021 166 1058 229
rect 1012 158 1058 166
rect 1060 158 1098 229
rect 1100 294 1105 302
rect 1100 238 1102 294
rect 1100 229 1105 238
rect 1107 229 1170 302
rect 1172 270 1210 302
rect 1172 229 1219 270
rect 1100 158 1140 229
rect 1142 158 1205 229
rect 1210 190 1219 229
rect 98 77 138 149
rect 140 77 203 149
rect 204 141 293 149
rect 213 85 293 141
rect 204 77 293 85
rect 295 77 398 149
rect 400 77 543 149
rect 545 77 648 149
rect 650 77 793 149
rect 795 77 898 149
rect 900 77 1043 149
rect 1045 122 1148 149
rect 1150 122 1213 149
rect 1045 120 1213 122
rect 1045 77 1148 120
rect 1150 77 1213 120
rect 5 75 101 77
rect 103 75 246 77
rect 248 75 351 77
rect 353 75 496 77
rect 498 75 601 77
rect 603 75 746 77
rect 748 75 851 77
rect 853 75 916 77
rect 917 75 1012 77
rect 5 5 85 75
rect 87 22 190 75
rect 87 13 100 22
rect 102 13 190 22
rect 87 5 190 13
rect 192 5 335 75
rect 337 5 440 75
rect 442 5 585 75
rect 587 5 690 75
rect 692 5 835 75
rect 837 71 1012 75
rect 837 34 940 71
rect 942 34 1005 71
rect 837 32 1005 34
rect 837 5 940 32
rect 942 5 1005 32
<< nwell >>
rect -5 306 211 386
rect 477 308 898 388
rect 477 269 1219 270
rect -5 268 1219 269
rect -6 190 1219 268
rect -6 117 94 118
rect -6 37 1218 117
<< pwell >>
rect -5 386 211 423
rect 477 388 898 425
rect 477 307 898 308
rect 211 306 1219 307
rect -5 270 1219 306
rect -5 269 477 270
rect -6 151 1219 190
rect -6 118 1218 151
rect 94 117 1218 118
rect -6 1 1219 37
rect -6 0 345 1
rect 561 0 1219 1
<< poly >>
rect 21 405 23 410
rect 28 405 30 410
rect 41 403 43 407
rect 61 405 63 410
rect 68 405 70 410
rect 126 414 151 416
rect 109 409 111 414
rect 116 409 118 414
rect 81 403 83 407
rect 126 406 128 414
rect 136 406 138 410
rect 149 406 151 414
rect 149 404 154 406
rect 173 405 175 410
rect 180 405 182 410
rect 503 407 505 412
rect 510 407 512 412
rect 152 401 154 404
rect 21 381 23 394
rect 28 389 30 394
rect 41 389 43 394
rect 27 387 33 389
rect 27 385 29 387
rect 31 385 33 387
rect 27 383 33 385
rect 37 387 43 389
rect 37 385 39 387
rect 41 385 43 387
rect 37 383 43 385
rect 17 379 23 381
rect 17 377 19 379
rect 21 377 23 379
rect 17 375 23 377
rect 21 372 23 375
rect 31 372 33 383
rect 41 379 43 383
rect 61 381 63 394
rect 68 389 70 394
rect 81 389 83 394
rect 67 387 73 389
rect 67 385 69 387
rect 71 385 73 387
rect 67 383 73 385
rect 77 387 83 389
rect 109 388 111 397
rect 116 394 118 397
rect 116 392 120 394
rect 126 393 128 397
rect 136 394 138 397
rect 118 389 120 392
rect 136 392 145 394
rect 193 403 195 407
rect 523 405 525 409
rect 543 407 545 412
rect 550 407 552 412
rect 608 416 633 418
rect 591 411 593 416
rect 598 411 600 416
rect 563 405 565 409
rect 608 408 610 416
rect 618 408 620 412
rect 631 408 633 416
rect 631 406 636 408
rect 655 407 657 412
rect 662 407 664 412
rect 634 403 636 406
rect 136 390 141 392
rect 143 390 145 392
rect 77 385 79 387
rect 81 385 83 387
rect 77 383 83 385
rect 57 379 63 381
rect 57 377 59 379
rect 61 377 63 379
rect 57 375 63 377
rect 61 372 63 375
rect 71 372 73 383
rect 81 379 83 383
rect 108 386 114 388
rect 108 384 110 386
rect 112 384 114 386
rect 108 382 114 384
rect 118 387 124 389
rect 118 385 120 387
rect 122 385 124 387
rect 118 383 124 385
rect 136 388 145 390
rect 136 384 138 388
rect 152 384 154 392
rect 108 379 110 382
rect 118 379 120 383
rect 128 382 138 384
rect 144 382 157 384
rect 128 379 130 382
rect 144 379 146 382
rect 155 381 157 382
rect 173 381 175 394
rect 180 389 182 394
rect 193 389 195 394
rect 179 387 185 389
rect 179 385 181 387
rect 183 385 185 387
rect 179 383 185 385
rect 189 387 195 389
rect 189 385 191 387
rect 193 385 195 387
rect 189 383 195 385
rect 503 383 505 396
rect 510 391 512 396
rect 523 391 525 396
rect 509 389 515 391
rect 509 387 511 389
rect 513 387 515 389
rect 509 385 515 387
rect 519 389 525 391
rect 519 387 521 389
rect 523 387 525 389
rect 519 385 525 387
rect 155 379 161 381
rect 21 354 23 359
rect 31 354 33 359
rect 41 357 43 361
rect 61 354 63 359
rect 71 354 73 359
rect 81 357 83 361
rect 118 357 120 361
rect 128 357 130 361
rect 108 348 110 352
rect 155 377 157 379
rect 159 377 161 379
rect 155 375 161 377
rect 169 379 175 381
rect 169 377 171 379
rect 173 377 175 379
rect 169 375 175 377
rect 173 372 175 375
rect 183 372 185 383
rect 193 379 195 383
rect 499 381 505 383
rect 499 379 501 381
rect 503 379 505 381
rect 499 377 505 379
rect 503 374 505 377
rect 513 374 515 385
rect 523 381 525 385
rect 543 383 545 396
rect 550 391 552 396
rect 563 391 565 396
rect 549 389 555 391
rect 549 387 551 389
rect 553 387 555 389
rect 549 385 555 387
rect 559 389 565 391
rect 591 390 593 399
rect 598 396 600 399
rect 598 394 602 396
rect 608 395 610 399
rect 618 396 620 399
rect 600 391 602 394
rect 618 394 627 396
rect 675 405 677 409
rect 708 407 710 412
rect 715 407 717 412
rect 728 405 730 409
rect 748 407 750 412
rect 755 407 757 412
rect 813 416 838 418
rect 796 411 798 416
rect 803 411 805 416
rect 768 405 770 409
rect 813 408 815 416
rect 823 408 825 412
rect 836 408 838 416
rect 836 406 841 408
rect 860 407 862 412
rect 867 407 869 412
rect 839 403 841 406
rect 618 392 623 394
rect 625 392 627 394
rect 559 387 561 389
rect 563 387 565 389
rect 559 385 565 387
rect 539 381 545 383
rect 539 379 541 381
rect 543 379 545 381
rect 539 377 545 379
rect 543 374 545 377
rect 553 374 555 385
rect 563 381 565 385
rect 590 388 596 390
rect 590 386 592 388
rect 594 386 596 388
rect 590 384 596 386
rect 600 389 606 391
rect 600 387 602 389
rect 604 387 606 389
rect 600 385 606 387
rect 618 390 627 392
rect 618 386 620 390
rect 634 386 636 394
rect 590 381 592 384
rect 600 381 602 385
rect 610 384 620 386
rect 626 384 639 386
rect 610 381 612 384
rect 626 381 628 384
rect 637 383 639 384
rect 655 383 657 396
rect 662 391 664 396
rect 675 391 677 396
rect 661 389 667 391
rect 661 387 663 389
rect 665 387 667 389
rect 661 385 667 387
rect 671 389 677 391
rect 671 387 673 389
rect 675 387 677 389
rect 671 385 677 387
rect 637 381 643 383
rect 173 354 175 359
rect 183 354 185 359
rect 193 357 195 361
rect 503 356 505 361
rect 513 356 515 361
rect 523 359 525 363
rect 543 356 545 361
rect 553 356 555 361
rect 563 359 565 363
rect 144 348 146 352
rect 600 359 602 363
rect 610 359 612 363
rect 590 350 592 354
rect 637 379 639 381
rect 641 379 643 381
rect 637 377 643 379
rect 651 381 657 383
rect 651 379 653 381
rect 655 379 657 381
rect 651 377 657 379
rect 655 374 657 377
rect 665 374 667 385
rect 675 381 677 385
rect 708 383 710 396
rect 715 391 717 396
rect 728 391 730 396
rect 714 389 720 391
rect 714 387 716 389
rect 718 387 720 389
rect 714 385 720 387
rect 724 389 730 391
rect 724 387 726 389
rect 728 387 730 389
rect 724 385 730 387
rect 704 381 710 383
rect 704 379 706 381
rect 708 379 710 381
rect 704 377 710 379
rect 708 374 710 377
rect 718 374 720 385
rect 728 381 730 385
rect 748 383 750 396
rect 755 391 757 396
rect 768 391 770 396
rect 754 389 760 391
rect 754 387 756 389
rect 758 387 760 389
rect 754 385 760 387
rect 764 389 770 391
rect 796 390 798 399
rect 803 396 805 399
rect 803 394 807 396
rect 813 395 815 399
rect 823 396 825 399
rect 805 391 807 394
rect 823 394 832 396
rect 880 405 882 409
rect 823 392 828 394
rect 830 392 832 394
rect 764 387 766 389
rect 768 387 770 389
rect 764 385 770 387
rect 744 381 750 383
rect 655 356 657 361
rect 665 356 667 361
rect 675 359 677 363
rect 744 379 746 381
rect 748 379 750 381
rect 744 377 750 379
rect 748 374 750 377
rect 758 374 760 385
rect 768 381 770 385
rect 795 388 801 390
rect 795 386 797 388
rect 799 386 801 388
rect 795 384 801 386
rect 805 389 811 391
rect 805 387 807 389
rect 809 387 811 389
rect 805 385 811 387
rect 823 390 832 392
rect 823 386 825 390
rect 839 386 841 394
rect 795 381 797 384
rect 805 381 807 385
rect 815 384 825 386
rect 831 384 844 386
rect 815 381 817 384
rect 831 381 833 384
rect 842 383 844 384
rect 860 383 862 396
rect 867 391 869 396
rect 880 391 882 396
rect 866 389 872 391
rect 866 387 868 389
rect 870 387 872 389
rect 866 385 872 387
rect 876 389 882 391
rect 876 387 878 389
rect 880 387 882 389
rect 876 385 882 387
rect 842 381 848 383
rect 708 356 710 361
rect 718 356 720 361
rect 728 359 730 363
rect 626 350 628 354
rect 748 356 750 361
rect 758 356 760 361
rect 768 359 770 363
rect 805 359 807 363
rect 815 359 817 363
rect 795 350 797 354
rect 842 379 844 381
rect 846 379 848 381
rect 842 377 848 379
rect 856 381 862 383
rect 856 379 858 381
rect 860 379 862 381
rect 856 377 862 379
rect 860 374 862 377
rect 870 374 872 385
rect 880 381 882 385
rect 860 356 862 361
rect 870 356 872 361
rect 880 359 882 363
rect 831 350 833 354
rect 21 331 23 335
rect 31 333 33 338
rect 41 333 43 338
rect 61 333 63 338
rect 71 333 73 338
rect 150 340 152 344
rect 81 331 83 335
rect 101 331 103 335
rect 111 333 113 338
rect 121 333 123 338
rect 21 309 23 313
rect 31 309 33 320
rect 41 317 43 320
rect 61 317 63 320
rect 41 315 47 317
rect 41 313 43 315
rect 45 313 47 315
rect 41 311 47 313
rect 57 315 63 317
rect 57 313 59 315
rect 61 313 63 315
rect 57 311 63 313
rect 21 307 27 309
rect 21 305 23 307
rect 25 305 27 307
rect 21 303 27 305
rect 31 307 37 309
rect 31 305 33 307
rect 35 305 37 307
rect 31 303 37 305
rect 21 298 23 303
rect 34 298 36 303
rect 41 298 43 311
rect 61 298 63 311
rect 71 309 73 320
rect 81 309 83 313
rect 67 307 73 309
rect 67 305 69 307
rect 71 305 73 307
rect 67 303 73 305
rect 77 307 83 309
rect 77 305 79 307
rect 81 305 83 307
rect 77 303 83 305
rect 68 298 70 303
rect 81 298 83 303
rect 101 309 103 313
rect 111 309 113 320
rect 121 317 123 320
rect 121 315 127 317
rect 121 313 123 315
rect 125 313 127 315
rect 121 311 127 313
rect 135 315 141 317
rect 135 313 137 315
rect 139 313 141 315
rect 186 340 188 344
rect 166 331 168 335
rect 176 331 178 335
rect 503 333 505 337
rect 513 335 515 340
rect 523 335 525 340
rect 543 335 545 340
rect 553 335 555 340
rect 632 342 634 346
rect 563 333 565 337
rect 583 333 585 337
rect 593 335 595 340
rect 603 335 605 340
rect 135 311 141 313
rect 101 307 107 309
rect 101 305 103 307
rect 105 305 107 307
rect 101 303 107 305
rect 111 307 117 309
rect 111 305 113 307
rect 115 305 117 307
rect 111 303 117 305
rect 101 298 103 303
rect 114 298 116 303
rect 121 298 123 311
rect 139 310 141 311
rect 150 310 152 313
rect 166 310 168 313
rect 139 308 152 310
rect 158 308 168 310
rect 176 309 178 313
rect 186 310 188 313
rect 142 300 144 308
rect 158 304 160 308
rect 151 302 160 304
rect 172 307 178 309
rect 172 305 174 307
rect 176 305 178 307
rect 172 303 178 305
rect 182 308 188 310
rect 182 306 184 308
rect 186 306 188 308
rect 182 304 188 306
rect 503 311 505 315
rect 513 311 515 322
rect 523 319 525 322
rect 543 319 545 322
rect 523 317 529 319
rect 523 315 525 317
rect 527 315 529 317
rect 523 313 529 315
rect 539 317 545 319
rect 539 315 541 317
rect 543 315 545 317
rect 539 313 545 315
rect 503 309 509 311
rect 503 307 505 309
rect 507 307 509 309
rect 503 305 509 307
rect 513 309 519 311
rect 513 307 515 309
rect 517 307 519 309
rect 513 305 519 307
rect 151 300 153 302
rect 155 300 160 302
rect 21 285 23 289
rect 34 282 36 287
rect 41 282 43 287
rect 61 282 63 287
rect 68 282 70 287
rect 81 285 83 289
rect 101 285 103 289
rect 151 298 160 300
rect 176 300 178 303
rect 158 295 160 298
rect 168 295 170 299
rect 176 298 180 300
rect 178 295 180 298
rect 185 295 187 304
rect 503 300 505 305
rect 516 300 518 305
rect 523 300 525 313
rect 543 300 545 313
rect 553 311 555 322
rect 563 311 565 315
rect 549 309 555 311
rect 549 307 551 309
rect 553 307 555 309
rect 549 305 555 307
rect 559 309 565 311
rect 559 307 561 309
rect 563 307 565 309
rect 559 305 565 307
rect 550 300 552 305
rect 563 300 565 305
rect 583 311 585 315
rect 593 311 595 322
rect 603 319 605 322
rect 603 317 609 319
rect 603 315 605 317
rect 607 315 609 317
rect 603 313 609 315
rect 617 317 623 319
rect 617 315 619 317
rect 621 315 623 317
rect 668 342 670 346
rect 648 333 650 337
rect 658 333 660 337
rect 708 333 710 337
rect 718 335 720 340
rect 728 335 730 340
rect 748 335 750 340
rect 758 335 760 340
rect 837 342 839 346
rect 768 333 770 337
rect 788 333 790 337
rect 798 335 800 340
rect 808 335 810 340
rect 617 313 623 315
rect 583 309 589 311
rect 583 307 585 309
rect 587 307 589 309
rect 583 305 589 307
rect 593 309 599 311
rect 593 307 595 309
rect 597 307 599 309
rect 593 305 599 307
rect 583 300 585 305
rect 596 300 598 305
rect 603 300 605 313
rect 621 312 623 313
rect 632 312 634 315
rect 648 312 650 315
rect 621 310 634 312
rect 640 310 650 312
rect 658 311 660 315
rect 668 312 670 315
rect 624 302 626 310
rect 640 306 642 310
rect 633 304 642 306
rect 654 309 660 311
rect 654 307 656 309
rect 658 307 660 309
rect 654 305 660 307
rect 664 310 670 312
rect 664 308 666 310
rect 668 308 670 310
rect 664 306 670 308
rect 708 311 710 315
rect 718 311 720 322
rect 728 319 730 322
rect 748 319 750 322
rect 728 317 734 319
rect 728 315 730 317
rect 732 315 734 317
rect 728 313 734 315
rect 744 317 750 319
rect 744 315 746 317
rect 748 315 750 317
rect 744 313 750 315
rect 708 309 714 311
rect 708 307 710 309
rect 712 307 714 309
rect 633 302 635 304
rect 637 302 642 304
rect 142 288 144 291
rect 114 282 116 287
rect 121 282 123 287
rect 142 286 147 288
rect 145 278 147 286
rect 158 282 160 286
rect 168 278 170 286
rect 503 287 505 291
rect 178 278 180 283
rect 185 278 187 283
rect 516 284 518 289
rect 523 284 525 289
rect 543 284 545 289
rect 550 284 552 289
rect 563 287 565 291
rect 583 287 585 291
rect 633 300 642 302
rect 658 302 660 305
rect 640 297 642 300
rect 650 297 652 301
rect 658 300 662 302
rect 660 297 662 300
rect 667 297 669 306
rect 708 305 714 307
rect 718 309 724 311
rect 718 307 720 309
rect 722 307 724 309
rect 718 305 724 307
rect 708 300 710 305
rect 721 300 723 305
rect 728 300 730 313
rect 748 300 750 313
rect 758 311 760 322
rect 768 311 770 315
rect 754 309 760 311
rect 754 307 756 309
rect 758 307 760 309
rect 754 305 760 307
rect 764 309 770 311
rect 764 307 766 309
rect 768 307 770 309
rect 764 305 770 307
rect 755 300 757 305
rect 768 300 770 305
rect 788 311 790 315
rect 798 311 800 322
rect 808 319 810 322
rect 808 317 814 319
rect 808 315 810 317
rect 812 315 814 317
rect 808 313 814 315
rect 822 317 828 319
rect 822 315 824 317
rect 826 315 828 317
rect 873 342 875 346
rect 853 333 855 337
rect 863 333 865 337
rect 822 313 828 315
rect 788 309 794 311
rect 788 307 790 309
rect 792 307 794 309
rect 788 305 794 307
rect 798 309 804 311
rect 798 307 800 309
rect 802 307 804 309
rect 798 305 804 307
rect 788 300 790 305
rect 801 300 803 305
rect 808 300 810 313
rect 826 312 828 313
rect 837 312 839 315
rect 853 312 855 315
rect 826 310 839 312
rect 845 310 855 312
rect 863 311 865 315
rect 873 312 875 315
rect 829 302 831 310
rect 845 306 847 310
rect 838 304 847 306
rect 859 309 865 311
rect 859 307 861 309
rect 863 307 865 309
rect 859 305 865 307
rect 869 310 875 312
rect 869 308 871 310
rect 873 308 875 310
rect 869 306 875 308
rect 838 302 840 304
rect 842 302 847 304
rect 624 290 626 293
rect 596 284 598 289
rect 603 284 605 289
rect 624 288 629 290
rect 627 280 629 288
rect 640 284 642 288
rect 650 280 652 288
rect 708 287 710 291
rect 660 280 662 285
rect 667 280 669 285
rect 145 276 170 278
rect 627 278 652 280
rect 721 284 723 289
rect 728 284 730 289
rect 748 284 750 289
rect 755 284 757 289
rect 768 287 770 291
rect 788 287 790 291
rect 838 300 847 302
rect 863 302 865 305
rect 845 297 847 300
rect 855 297 857 301
rect 863 300 867 302
rect 865 297 867 300
rect 872 297 874 306
rect 829 290 831 293
rect 801 284 803 289
rect 808 284 810 289
rect 829 288 834 290
rect 832 280 834 288
rect 845 284 847 288
rect 855 280 857 288
rect 1029 289 1031 294
rect 1036 289 1038 294
rect 865 280 867 285
rect 872 280 874 285
rect 832 278 857 280
rect 1049 287 1051 291
rect 1069 289 1071 294
rect 1076 289 1078 294
rect 1134 298 1159 300
rect 1117 293 1119 298
rect 1124 293 1126 298
rect 1089 287 1091 291
rect 1134 290 1136 298
rect 1144 290 1146 294
rect 1157 290 1159 298
rect 1157 288 1162 290
rect 1181 289 1183 294
rect 1188 289 1190 294
rect 1160 285 1162 288
rect 1029 265 1031 278
rect 1036 273 1038 278
rect 1049 273 1051 278
rect 1035 271 1041 273
rect 1035 269 1037 271
rect 1039 269 1041 271
rect 1035 267 1041 269
rect 1045 271 1051 273
rect 1045 269 1047 271
rect 1049 269 1051 271
rect 1045 267 1051 269
rect 1025 263 1031 265
rect 1025 261 1027 263
rect 1029 261 1031 263
rect 1025 259 1031 261
rect 1029 256 1031 259
rect 1039 256 1041 267
rect 1049 263 1051 267
rect 1069 265 1071 278
rect 1076 273 1078 278
rect 1089 273 1091 278
rect 1075 271 1081 273
rect 1075 269 1077 271
rect 1079 269 1081 271
rect 1075 267 1081 269
rect 1085 271 1091 273
rect 1117 272 1119 281
rect 1124 278 1126 281
rect 1124 276 1128 278
rect 1134 277 1136 281
rect 1144 278 1146 281
rect 1126 273 1128 276
rect 1144 276 1153 278
rect 1201 287 1203 291
rect 1144 274 1149 276
rect 1151 274 1153 276
rect 1085 269 1087 271
rect 1089 269 1091 271
rect 1085 267 1091 269
rect 1065 263 1071 265
rect 1065 261 1067 263
rect 1069 261 1071 263
rect 1065 259 1071 261
rect 1069 256 1071 259
rect 1079 256 1081 267
rect 1089 263 1091 267
rect 1116 270 1122 272
rect 1116 268 1118 270
rect 1120 268 1122 270
rect 1116 266 1122 268
rect 1126 271 1132 273
rect 1126 269 1128 271
rect 1130 269 1132 271
rect 1126 267 1132 269
rect 1144 272 1153 274
rect 1144 268 1146 272
rect 1160 268 1162 276
rect 1116 263 1118 266
rect 1126 263 1128 267
rect 1136 266 1146 268
rect 1152 266 1165 268
rect 1136 263 1138 266
rect 1152 263 1154 266
rect 1163 265 1165 266
rect 1181 265 1183 278
rect 1188 273 1190 278
rect 1201 273 1203 278
rect 1187 271 1193 273
rect 1187 269 1189 271
rect 1191 269 1193 271
rect 1187 267 1193 269
rect 1197 271 1203 273
rect 1197 269 1199 271
rect 1201 269 1203 271
rect 1197 267 1203 269
rect 1163 263 1169 265
rect 1029 238 1031 243
rect 1039 238 1041 243
rect 1049 241 1051 245
rect 1069 238 1071 243
rect 1079 238 1081 243
rect 1089 241 1091 245
rect 1126 241 1128 245
rect 1136 241 1138 245
rect 1116 232 1118 236
rect 1163 261 1165 263
rect 1167 261 1169 263
rect 1163 259 1169 261
rect 1177 263 1183 265
rect 1177 261 1179 263
rect 1181 261 1183 263
rect 1177 259 1183 261
rect 1181 256 1183 259
rect 1191 256 1193 267
rect 1201 263 1203 267
rect 1181 238 1183 243
rect 1191 238 1193 243
rect 1201 241 1203 245
rect 1152 232 1154 236
rect 21 224 23 228
rect 28 224 30 228
rect 8 214 10 219
rect 97 224 99 228
rect 48 215 50 219
rect 58 217 60 222
rect 68 217 70 222
rect 8 193 10 196
rect 21 193 23 203
rect 28 200 30 203
rect 28 198 34 200
rect 28 196 30 198
rect 32 196 34 198
rect 28 194 34 196
rect 8 191 14 193
rect 8 189 10 191
rect 12 189 14 191
rect 8 187 14 189
rect 18 191 24 193
rect 18 189 20 191
rect 22 189 24 191
rect 18 187 24 189
rect 8 184 10 187
rect 18 184 20 187
rect 28 184 30 194
rect 48 193 50 197
rect 58 193 60 204
rect 68 201 70 204
rect 68 199 74 201
rect 68 197 70 199
rect 72 197 74 199
rect 68 195 74 197
rect 82 199 88 201
rect 82 197 84 199
rect 86 197 88 199
rect 133 224 135 228
rect 113 215 115 219
rect 123 215 125 219
rect 202 224 204 228
rect 153 215 155 219
rect 163 217 165 222
rect 173 217 175 222
rect 82 195 88 197
rect 48 191 54 193
rect 48 189 50 191
rect 52 189 54 191
rect 48 187 54 189
rect 58 191 64 193
rect 58 189 60 191
rect 62 189 64 191
rect 58 187 64 189
rect 48 182 50 187
rect 61 182 63 187
rect 68 182 70 195
rect 86 194 88 195
rect 97 194 99 197
rect 113 194 115 197
rect 86 192 99 194
rect 105 192 115 194
rect 123 193 125 197
rect 133 194 135 197
rect 89 184 91 192
rect 105 188 107 192
rect 98 186 107 188
rect 119 191 125 193
rect 119 189 121 191
rect 123 189 125 191
rect 119 187 125 189
rect 129 192 135 194
rect 129 190 131 192
rect 133 190 135 192
rect 129 188 135 190
rect 153 193 155 197
rect 163 193 165 204
rect 173 201 175 204
rect 173 199 179 201
rect 173 197 175 199
rect 177 197 179 199
rect 173 195 179 197
rect 187 199 193 201
rect 187 197 189 199
rect 191 197 193 199
rect 238 224 240 228
rect 218 215 220 219
rect 228 215 230 219
rect 271 224 273 228
rect 278 224 280 228
rect 258 214 260 219
rect 187 195 193 197
rect 153 191 159 193
rect 153 189 155 191
rect 157 189 159 191
rect 98 184 100 186
rect 102 184 107 186
rect 8 170 10 175
rect 18 173 20 178
rect 28 173 30 178
rect 48 169 50 173
rect 98 182 107 184
rect 123 184 125 187
rect 105 179 107 182
rect 115 179 117 183
rect 123 182 127 184
rect 125 179 127 182
rect 132 179 134 188
rect 153 187 159 189
rect 163 191 169 193
rect 163 189 165 191
rect 167 189 169 191
rect 163 187 169 189
rect 153 182 155 187
rect 166 182 168 187
rect 173 182 175 195
rect 191 194 193 195
rect 202 194 204 197
rect 218 194 220 197
rect 191 192 204 194
rect 210 192 220 194
rect 228 193 230 197
rect 238 194 240 197
rect 347 224 349 228
rect 298 215 300 219
rect 308 217 310 222
rect 318 217 320 222
rect 194 184 196 192
rect 210 188 212 192
rect 203 186 212 188
rect 224 191 230 193
rect 224 189 226 191
rect 228 189 230 191
rect 224 187 230 189
rect 234 192 240 194
rect 234 190 236 192
rect 238 190 240 192
rect 234 188 240 190
rect 258 193 260 196
rect 271 193 273 203
rect 278 200 280 203
rect 278 198 284 200
rect 278 196 280 198
rect 282 196 284 198
rect 278 194 284 196
rect 258 191 264 193
rect 258 189 260 191
rect 262 189 264 191
rect 203 184 205 186
rect 207 184 212 186
rect 89 172 91 175
rect 61 166 63 171
rect 68 166 70 171
rect 89 170 94 172
rect 92 162 94 170
rect 105 166 107 170
rect 115 162 117 170
rect 153 169 155 173
rect 203 182 212 184
rect 228 184 230 187
rect 210 179 212 182
rect 220 179 222 183
rect 228 182 232 184
rect 230 179 232 182
rect 237 179 239 188
rect 258 187 264 189
rect 268 191 274 193
rect 268 189 270 191
rect 272 189 274 191
rect 268 187 274 189
rect 258 184 260 187
rect 268 184 270 187
rect 278 184 280 194
rect 298 193 300 197
rect 308 193 310 204
rect 318 201 320 204
rect 318 199 324 201
rect 318 197 320 199
rect 322 197 324 199
rect 318 195 324 197
rect 332 199 338 201
rect 332 197 334 199
rect 336 197 338 199
rect 383 224 385 228
rect 363 215 365 219
rect 373 215 375 219
rect 452 224 454 228
rect 403 215 405 219
rect 413 217 415 222
rect 423 217 425 222
rect 332 195 338 197
rect 298 191 304 193
rect 298 189 300 191
rect 302 189 304 191
rect 298 187 304 189
rect 308 191 314 193
rect 308 189 310 191
rect 312 189 314 191
rect 308 187 314 189
rect 194 172 196 175
rect 125 162 127 167
rect 132 162 134 167
rect 92 160 117 162
rect 166 166 168 171
rect 173 166 175 171
rect 194 170 199 172
rect 197 162 199 170
rect 210 166 212 170
rect 220 162 222 170
rect 298 182 300 187
rect 311 182 313 187
rect 318 182 320 195
rect 336 194 338 195
rect 347 194 349 197
rect 363 194 365 197
rect 336 192 349 194
rect 355 192 365 194
rect 373 193 375 197
rect 383 194 385 197
rect 339 184 341 192
rect 355 188 357 192
rect 348 186 357 188
rect 369 191 375 193
rect 369 189 371 191
rect 373 189 375 191
rect 369 187 375 189
rect 379 192 385 194
rect 379 190 381 192
rect 383 190 385 192
rect 379 188 385 190
rect 403 193 405 197
rect 413 193 415 204
rect 423 201 425 204
rect 423 199 429 201
rect 423 197 425 199
rect 427 197 429 199
rect 423 195 429 197
rect 437 199 443 201
rect 437 197 439 199
rect 441 197 443 199
rect 488 224 490 228
rect 468 215 470 219
rect 478 215 480 219
rect 521 224 523 228
rect 528 224 530 228
rect 508 214 510 219
rect 437 195 443 197
rect 403 191 409 193
rect 403 189 405 191
rect 407 189 409 191
rect 348 184 350 186
rect 352 184 357 186
rect 258 170 260 175
rect 268 173 270 178
rect 278 173 280 178
rect 230 162 232 167
rect 237 162 239 167
rect 197 160 222 162
rect 298 169 300 173
rect 348 182 357 184
rect 373 184 375 187
rect 355 179 357 182
rect 365 179 367 183
rect 373 182 377 184
rect 375 179 377 182
rect 382 179 384 188
rect 403 187 409 189
rect 413 191 419 193
rect 413 189 415 191
rect 417 189 419 191
rect 413 187 419 189
rect 403 182 405 187
rect 416 182 418 187
rect 423 182 425 195
rect 441 194 443 195
rect 452 194 454 197
rect 468 194 470 197
rect 441 192 454 194
rect 460 192 470 194
rect 478 193 480 197
rect 488 194 490 197
rect 597 224 599 228
rect 548 215 550 219
rect 558 217 560 222
rect 568 217 570 222
rect 444 184 446 192
rect 460 188 462 192
rect 453 186 462 188
rect 474 191 480 193
rect 474 189 476 191
rect 478 189 480 191
rect 474 187 480 189
rect 484 192 490 194
rect 484 190 486 192
rect 488 190 490 192
rect 484 188 490 190
rect 508 193 510 196
rect 521 193 523 203
rect 528 200 530 203
rect 528 198 534 200
rect 528 196 530 198
rect 532 196 534 198
rect 528 194 534 196
rect 508 191 514 193
rect 508 189 510 191
rect 512 189 514 191
rect 453 184 455 186
rect 457 184 462 186
rect 339 172 341 175
rect 311 166 313 171
rect 318 166 320 171
rect 339 170 344 172
rect 342 162 344 170
rect 355 166 357 170
rect 365 162 367 170
rect 403 169 405 173
rect 453 182 462 184
rect 478 184 480 187
rect 460 179 462 182
rect 470 179 472 183
rect 478 182 482 184
rect 480 179 482 182
rect 487 179 489 188
rect 508 187 514 189
rect 518 191 524 193
rect 518 189 520 191
rect 522 189 524 191
rect 518 187 524 189
rect 508 184 510 187
rect 518 184 520 187
rect 528 184 530 194
rect 548 193 550 197
rect 558 193 560 204
rect 568 201 570 204
rect 568 199 574 201
rect 568 197 570 199
rect 572 197 574 199
rect 568 195 574 197
rect 582 199 588 201
rect 582 197 584 199
rect 586 197 588 199
rect 633 224 635 228
rect 613 215 615 219
rect 623 215 625 219
rect 702 224 704 228
rect 653 215 655 219
rect 663 217 665 222
rect 673 217 675 222
rect 582 195 588 197
rect 548 191 554 193
rect 548 189 550 191
rect 552 189 554 191
rect 548 187 554 189
rect 558 191 564 193
rect 558 189 560 191
rect 562 189 564 191
rect 558 187 564 189
rect 444 172 446 175
rect 375 162 377 167
rect 382 162 384 167
rect 342 160 367 162
rect 416 166 418 171
rect 423 166 425 171
rect 444 170 449 172
rect 447 162 449 170
rect 460 166 462 170
rect 470 162 472 170
rect 548 182 550 187
rect 561 182 563 187
rect 568 182 570 195
rect 586 194 588 195
rect 597 194 599 197
rect 613 194 615 197
rect 586 192 599 194
rect 605 192 615 194
rect 623 193 625 197
rect 633 194 635 197
rect 589 184 591 192
rect 605 188 607 192
rect 598 186 607 188
rect 619 191 625 193
rect 619 189 621 191
rect 623 189 625 191
rect 619 187 625 189
rect 629 192 635 194
rect 629 190 631 192
rect 633 190 635 192
rect 629 188 635 190
rect 653 193 655 197
rect 663 193 665 204
rect 673 201 675 204
rect 673 199 679 201
rect 673 197 675 199
rect 677 197 679 199
rect 673 195 679 197
rect 687 199 693 201
rect 687 197 689 199
rect 691 197 693 199
rect 738 224 740 228
rect 718 215 720 219
rect 728 215 730 219
rect 771 224 773 228
rect 778 224 780 228
rect 758 214 760 219
rect 687 195 693 197
rect 653 191 659 193
rect 653 189 655 191
rect 657 189 659 191
rect 598 184 600 186
rect 602 184 607 186
rect 508 170 510 175
rect 518 173 520 178
rect 528 173 530 178
rect 480 162 482 167
rect 487 162 489 167
rect 447 160 472 162
rect 548 169 550 173
rect 598 182 607 184
rect 623 184 625 187
rect 605 179 607 182
rect 615 179 617 183
rect 623 182 627 184
rect 625 179 627 182
rect 632 179 634 188
rect 653 187 659 189
rect 663 191 669 193
rect 663 189 665 191
rect 667 189 669 191
rect 663 187 669 189
rect 653 182 655 187
rect 666 182 668 187
rect 673 182 675 195
rect 691 194 693 195
rect 702 194 704 197
rect 718 194 720 197
rect 691 192 704 194
rect 710 192 720 194
rect 728 193 730 197
rect 738 194 740 197
rect 847 224 849 228
rect 798 215 800 219
rect 808 217 810 222
rect 818 217 820 222
rect 694 184 696 192
rect 710 188 712 192
rect 703 186 712 188
rect 724 191 730 193
rect 724 189 726 191
rect 728 189 730 191
rect 724 187 730 189
rect 734 192 740 194
rect 734 190 736 192
rect 738 190 740 192
rect 734 188 740 190
rect 758 193 760 196
rect 771 193 773 203
rect 778 200 780 203
rect 778 198 784 200
rect 778 196 780 198
rect 782 196 784 198
rect 778 194 784 196
rect 758 191 764 193
rect 758 189 760 191
rect 762 189 764 191
rect 703 184 705 186
rect 707 184 712 186
rect 589 172 591 175
rect 561 166 563 171
rect 568 166 570 171
rect 589 170 594 172
rect 592 162 594 170
rect 605 166 607 170
rect 615 162 617 170
rect 653 169 655 173
rect 703 182 712 184
rect 728 184 730 187
rect 710 179 712 182
rect 720 179 722 183
rect 728 182 732 184
rect 730 179 732 182
rect 737 179 739 188
rect 758 187 764 189
rect 768 191 774 193
rect 768 189 770 191
rect 772 189 774 191
rect 768 187 774 189
rect 758 184 760 187
rect 768 184 770 187
rect 778 184 780 194
rect 798 193 800 197
rect 808 193 810 204
rect 818 201 820 204
rect 818 199 824 201
rect 818 197 820 199
rect 822 197 824 199
rect 818 195 824 197
rect 832 199 838 201
rect 832 197 834 199
rect 836 197 838 199
rect 883 224 885 228
rect 863 215 865 219
rect 873 215 875 219
rect 952 224 954 228
rect 903 215 905 219
rect 913 217 915 222
rect 923 217 925 222
rect 832 195 838 197
rect 798 191 804 193
rect 798 189 800 191
rect 802 189 804 191
rect 798 187 804 189
rect 808 191 814 193
rect 808 189 810 191
rect 812 189 814 191
rect 808 187 814 189
rect 694 172 696 175
rect 625 162 627 167
rect 632 162 634 167
rect 592 160 617 162
rect 666 166 668 171
rect 673 166 675 171
rect 694 170 699 172
rect 697 162 699 170
rect 710 166 712 170
rect 720 162 722 170
rect 798 182 800 187
rect 811 182 813 187
rect 818 182 820 195
rect 836 194 838 195
rect 847 194 849 197
rect 863 194 865 197
rect 836 192 849 194
rect 855 192 865 194
rect 873 193 875 197
rect 883 194 885 197
rect 839 184 841 192
rect 855 188 857 192
rect 848 186 857 188
rect 869 191 875 193
rect 869 189 871 191
rect 873 189 875 191
rect 869 187 875 189
rect 879 192 885 194
rect 879 190 881 192
rect 883 190 885 192
rect 879 188 885 190
rect 903 193 905 197
rect 913 193 915 204
rect 923 201 925 204
rect 923 199 929 201
rect 923 197 925 199
rect 927 197 929 199
rect 923 195 929 197
rect 937 199 943 201
rect 937 197 939 199
rect 941 197 943 199
rect 988 224 990 228
rect 968 215 970 219
rect 978 215 980 219
rect 1029 215 1031 219
rect 1039 217 1041 222
rect 1049 217 1051 222
rect 1069 217 1071 222
rect 1079 217 1081 222
rect 1158 224 1160 228
rect 1089 215 1091 219
rect 1109 215 1111 219
rect 1119 217 1121 222
rect 1129 217 1131 222
rect 937 195 943 197
rect 903 191 909 193
rect 903 189 905 191
rect 907 189 909 191
rect 848 184 850 186
rect 852 184 857 186
rect 758 170 760 175
rect 768 173 770 178
rect 778 173 780 178
rect 730 162 732 167
rect 737 162 739 167
rect 697 160 722 162
rect 798 169 800 173
rect 848 182 857 184
rect 873 184 875 187
rect 855 179 857 182
rect 865 179 867 183
rect 873 182 877 184
rect 875 179 877 182
rect 882 179 884 188
rect 903 187 909 189
rect 913 191 919 193
rect 913 189 915 191
rect 917 189 919 191
rect 913 187 919 189
rect 903 182 905 187
rect 916 182 918 187
rect 923 182 925 195
rect 941 194 943 195
rect 952 194 954 197
rect 968 194 970 197
rect 941 192 954 194
rect 960 192 970 194
rect 978 193 980 197
rect 988 194 990 197
rect 944 184 946 192
rect 960 188 962 192
rect 953 186 962 188
rect 974 191 980 193
rect 974 189 976 191
rect 978 189 980 191
rect 974 187 980 189
rect 984 192 990 194
rect 984 190 986 192
rect 988 190 990 192
rect 984 188 990 190
rect 1029 193 1031 197
rect 1039 193 1041 204
rect 1049 201 1051 204
rect 1069 201 1071 204
rect 1049 199 1055 201
rect 1049 197 1051 199
rect 1053 197 1055 199
rect 1049 195 1055 197
rect 1065 199 1071 201
rect 1065 197 1067 199
rect 1069 197 1071 199
rect 1065 195 1071 197
rect 1029 191 1035 193
rect 1029 189 1031 191
rect 1033 189 1035 191
rect 953 184 955 186
rect 957 184 962 186
rect 839 172 841 175
rect 811 166 813 171
rect 818 166 820 171
rect 839 170 844 172
rect 842 162 844 170
rect 855 166 857 170
rect 865 162 867 170
rect 903 169 905 173
rect 953 182 962 184
rect 978 184 980 187
rect 960 179 962 182
rect 970 179 972 183
rect 978 182 982 184
rect 980 179 982 182
rect 987 179 989 188
rect 1029 187 1035 189
rect 1039 191 1045 193
rect 1039 189 1041 191
rect 1043 189 1045 191
rect 1039 187 1045 189
rect 1029 182 1031 187
rect 1042 182 1044 187
rect 1049 182 1051 195
rect 1069 182 1071 195
rect 1079 193 1081 204
rect 1089 193 1091 197
rect 1075 191 1081 193
rect 1075 189 1077 191
rect 1079 189 1081 191
rect 1075 187 1081 189
rect 1085 191 1091 193
rect 1085 189 1087 191
rect 1089 189 1091 191
rect 1085 187 1091 189
rect 1076 182 1078 187
rect 1089 182 1091 187
rect 1109 193 1111 197
rect 1119 193 1121 204
rect 1129 201 1131 204
rect 1129 199 1135 201
rect 1129 197 1131 199
rect 1133 197 1135 199
rect 1129 195 1135 197
rect 1143 199 1149 201
rect 1143 197 1145 199
rect 1147 197 1149 199
rect 1194 224 1196 228
rect 1174 215 1176 219
rect 1184 215 1186 219
rect 1143 195 1149 197
rect 1109 191 1115 193
rect 1109 189 1111 191
rect 1113 189 1115 191
rect 1109 187 1115 189
rect 1119 191 1125 193
rect 1119 189 1121 191
rect 1123 189 1125 191
rect 1119 187 1125 189
rect 1109 182 1111 187
rect 1122 182 1124 187
rect 1129 182 1131 195
rect 1147 194 1149 195
rect 1158 194 1160 197
rect 1174 194 1176 197
rect 1147 192 1160 194
rect 1166 192 1176 194
rect 1184 193 1186 197
rect 1194 194 1196 197
rect 1150 184 1152 192
rect 1166 188 1168 192
rect 1159 186 1168 188
rect 1180 191 1186 193
rect 1180 189 1182 191
rect 1184 189 1186 191
rect 1180 187 1186 189
rect 1190 192 1196 194
rect 1190 190 1192 192
rect 1194 190 1196 192
rect 1190 188 1196 190
rect 1159 184 1161 186
rect 1163 184 1168 186
rect 944 172 946 175
rect 875 162 877 167
rect 882 162 884 167
rect 842 160 867 162
rect 916 166 918 171
rect 923 166 925 171
rect 944 170 949 172
rect 947 162 949 170
rect 960 166 962 170
rect 970 162 972 170
rect 1029 169 1031 173
rect 980 162 982 167
rect 987 162 989 167
rect 947 160 972 162
rect 1042 166 1044 171
rect 1049 166 1051 171
rect 1069 166 1071 171
rect 1076 166 1078 171
rect 1089 169 1091 173
rect 1109 169 1111 173
rect 1159 182 1168 184
rect 1184 184 1186 187
rect 1166 179 1168 182
rect 1176 179 1178 183
rect 1184 182 1188 184
rect 1186 179 1188 182
rect 1193 179 1195 188
rect 1150 172 1152 175
rect 1122 166 1124 171
rect 1129 166 1131 171
rect 1150 170 1155 172
rect 1153 162 1155 170
rect 1166 166 1168 170
rect 1176 162 1178 170
rect 1186 162 1188 167
rect 1193 162 1195 167
rect 1153 160 1178 162
rect 107 134 109 138
rect 120 136 122 141
rect 127 136 129 141
rect 151 145 176 147
rect 151 137 153 145
rect 164 137 166 141
rect 174 137 176 145
rect 184 140 186 145
rect 191 140 193 145
rect 148 135 153 137
rect 148 132 150 135
rect 107 120 109 125
rect 120 120 122 125
rect 107 118 113 120
rect 107 116 109 118
rect 111 116 113 118
rect 107 114 113 116
rect 117 118 123 120
rect 117 116 119 118
rect 121 116 123 118
rect 117 114 123 116
rect 107 110 109 114
rect 117 103 119 114
rect 127 112 129 125
rect 222 132 224 137
rect 164 125 166 128
rect 157 123 166 125
rect 174 124 176 128
rect 184 125 186 128
rect 148 115 150 123
rect 157 121 159 123
rect 161 121 166 123
rect 157 119 166 121
rect 182 123 186 125
rect 182 120 184 123
rect 164 115 166 119
rect 178 118 184 120
rect 191 119 193 128
rect 232 129 234 134
rect 242 129 244 134
rect 262 134 264 138
rect 275 136 277 141
rect 282 136 284 141
rect 306 145 331 147
rect 306 137 308 145
rect 319 137 321 141
rect 329 137 331 145
rect 339 140 341 145
rect 346 140 348 145
rect 303 135 308 137
rect 303 132 305 135
rect 222 120 224 123
rect 232 120 234 123
rect 178 116 180 118
rect 182 116 184 118
rect 145 113 158 115
rect 164 113 174 115
rect 178 114 184 116
rect 145 112 147 113
rect 127 110 133 112
rect 127 108 129 110
rect 131 108 133 110
rect 127 106 133 108
rect 141 110 147 112
rect 156 110 158 113
rect 172 110 174 113
rect 182 110 184 114
rect 188 117 194 119
rect 188 115 190 117
rect 192 115 194 117
rect 188 113 194 115
rect 192 110 194 113
rect 222 118 228 120
rect 222 116 224 118
rect 226 116 228 118
rect 222 114 228 116
rect 232 118 238 120
rect 232 116 234 118
rect 236 116 238 118
rect 232 114 238 116
rect 222 111 224 114
rect 141 108 143 110
rect 145 108 147 110
rect 141 106 147 108
rect 127 103 129 106
rect 107 88 109 92
rect 117 85 119 90
rect 127 85 129 90
rect 172 88 174 92
rect 182 88 184 92
rect 156 79 158 83
rect 235 104 237 114
rect 242 113 244 123
rect 262 120 264 125
rect 275 120 277 125
rect 262 118 268 120
rect 262 116 264 118
rect 266 116 268 118
rect 262 114 268 116
rect 272 118 278 120
rect 272 116 274 118
rect 276 116 278 118
rect 272 114 278 116
rect 242 111 248 113
rect 242 109 244 111
rect 246 109 248 111
rect 262 110 264 114
rect 242 107 248 109
rect 242 104 244 107
rect 222 88 224 93
rect 192 79 194 83
rect 272 103 274 114
rect 282 112 284 125
rect 367 134 369 138
rect 380 136 382 141
rect 387 136 389 141
rect 411 145 436 147
rect 411 137 413 145
rect 424 137 426 141
rect 434 137 436 145
rect 444 140 446 145
rect 451 140 453 145
rect 319 125 321 128
rect 312 123 321 125
rect 329 124 331 128
rect 339 125 341 128
rect 303 115 305 123
rect 312 121 314 123
rect 316 121 321 123
rect 312 119 321 121
rect 337 123 341 125
rect 337 120 339 123
rect 319 115 321 119
rect 333 118 339 120
rect 346 119 348 128
rect 408 135 413 137
rect 408 132 410 135
rect 367 120 369 125
rect 380 120 382 125
rect 333 116 335 118
rect 337 116 339 118
rect 300 113 313 115
rect 319 113 329 115
rect 333 114 339 116
rect 300 112 302 113
rect 282 110 288 112
rect 282 108 284 110
rect 286 108 288 110
rect 282 106 288 108
rect 296 110 302 112
rect 311 110 313 113
rect 327 110 329 113
rect 337 110 339 114
rect 343 117 349 119
rect 343 115 345 117
rect 347 115 349 117
rect 343 113 349 115
rect 347 110 349 113
rect 367 118 373 120
rect 367 116 369 118
rect 371 116 373 118
rect 367 114 373 116
rect 377 118 383 120
rect 377 116 379 118
rect 381 116 383 118
rect 377 114 383 116
rect 367 110 369 114
rect 296 108 298 110
rect 300 108 302 110
rect 296 106 302 108
rect 282 103 284 106
rect 262 88 264 92
rect 272 85 274 90
rect 282 85 284 90
rect 235 79 237 83
rect 242 79 244 83
rect 327 88 329 92
rect 337 88 339 92
rect 311 79 313 83
rect 377 103 379 114
rect 387 112 389 125
rect 472 132 474 137
rect 424 125 426 128
rect 417 123 426 125
rect 434 124 436 128
rect 444 125 446 128
rect 408 115 410 123
rect 417 121 419 123
rect 421 121 426 123
rect 417 119 426 121
rect 442 123 446 125
rect 442 120 444 123
rect 424 115 426 119
rect 438 118 444 120
rect 451 119 453 128
rect 482 129 484 134
rect 492 129 494 134
rect 512 134 514 138
rect 525 136 527 141
rect 532 136 534 141
rect 556 145 581 147
rect 556 137 558 145
rect 569 137 571 141
rect 579 137 581 145
rect 589 140 591 145
rect 596 140 598 145
rect 553 135 558 137
rect 553 132 555 135
rect 472 120 474 123
rect 482 120 484 123
rect 438 116 440 118
rect 442 116 444 118
rect 405 113 418 115
rect 424 113 434 115
rect 438 114 444 116
rect 405 112 407 113
rect 387 110 393 112
rect 387 108 389 110
rect 391 108 393 110
rect 387 106 393 108
rect 401 110 407 112
rect 416 110 418 113
rect 432 110 434 113
rect 442 110 444 114
rect 448 117 454 119
rect 448 115 450 117
rect 452 115 454 117
rect 448 113 454 115
rect 452 110 454 113
rect 472 118 478 120
rect 472 116 474 118
rect 476 116 478 118
rect 472 114 478 116
rect 482 118 488 120
rect 482 116 484 118
rect 486 116 488 118
rect 482 114 488 116
rect 472 111 474 114
rect 401 108 403 110
rect 405 108 407 110
rect 401 106 407 108
rect 387 103 389 106
rect 367 88 369 92
rect 377 85 379 90
rect 387 85 389 90
rect 347 79 349 83
rect 432 88 434 92
rect 442 88 444 92
rect 416 79 418 83
rect 485 104 487 114
rect 492 113 494 123
rect 512 120 514 125
rect 525 120 527 125
rect 512 118 518 120
rect 512 116 514 118
rect 516 116 518 118
rect 512 114 518 116
rect 522 118 528 120
rect 522 116 524 118
rect 526 116 528 118
rect 522 114 528 116
rect 492 111 498 113
rect 492 109 494 111
rect 496 109 498 111
rect 512 110 514 114
rect 492 107 498 109
rect 492 104 494 107
rect 472 88 474 93
rect 452 79 454 83
rect 522 103 524 114
rect 532 112 534 125
rect 617 134 619 138
rect 630 136 632 141
rect 637 136 639 141
rect 661 145 686 147
rect 661 137 663 145
rect 674 137 676 141
rect 684 137 686 145
rect 694 140 696 145
rect 701 140 703 145
rect 569 125 571 128
rect 562 123 571 125
rect 579 124 581 128
rect 589 125 591 128
rect 553 115 555 123
rect 562 121 564 123
rect 566 121 571 123
rect 562 119 571 121
rect 587 123 591 125
rect 587 120 589 123
rect 569 115 571 119
rect 583 118 589 120
rect 596 119 598 128
rect 658 135 663 137
rect 658 132 660 135
rect 617 120 619 125
rect 630 120 632 125
rect 583 116 585 118
rect 587 116 589 118
rect 550 113 563 115
rect 569 113 579 115
rect 583 114 589 116
rect 550 112 552 113
rect 532 110 538 112
rect 532 108 534 110
rect 536 108 538 110
rect 532 106 538 108
rect 546 110 552 112
rect 561 110 563 113
rect 577 110 579 113
rect 587 110 589 114
rect 593 117 599 119
rect 593 115 595 117
rect 597 115 599 117
rect 593 113 599 115
rect 597 110 599 113
rect 617 118 623 120
rect 617 116 619 118
rect 621 116 623 118
rect 617 114 623 116
rect 627 118 633 120
rect 627 116 629 118
rect 631 116 633 118
rect 627 114 633 116
rect 617 110 619 114
rect 546 108 548 110
rect 550 108 552 110
rect 546 106 552 108
rect 532 103 534 106
rect 512 88 514 92
rect 522 85 524 90
rect 532 85 534 90
rect 485 79 487 83
rect 492 79 494 83
rect 577 88 579 92
rect 587 88 589 92
rect 561 79 563 83
rect 627 103 629 114
rect 637 112 639 125
rect 722 132 724 137
rect 674 125 676 128
rect 667 123 676 125
rect 684 124 686 128
rect 694 125 696 128
rect 658 115 660 123
rect 667 121 669 123
rect 671 121 676 123
rect 667 119 676 121
rect 692 123 696 125
rect 692 120 694 123
rect 674 115 676 119
rect 688 118 694 120
rect 701 119 703 128
rect 732 129 734 134
rect 742 129 744 134
rect 762 134 764 138
rect 775 136 777 141
rect 782 136 784 141
rect 806 145 831 147
rect 806 137 808 145
rect 819 137 821 141
rect 829 137 831 145
rect 839 140 841 145
rect 846 140 848 145
rect 803 135 808 137
rect 803 132 805 135
rect 722 120 724 123
rect 732 120 734 123
rect 688 116 690 118
rect 692 116 694 118
rect 655 113 668 115
rect 674 113 684 115
rect 688 114 694 116
rect 655 112 657 113
rect 637 110 643 112
rect 637 108 639 110
rect 641 108 643 110
rect 637 106 643 108
rect 651 110 657 112
rect 666 110 668 113
rect 682 110 684 113
rect 692 110 694 114
rect 698 117 704 119
rect 698 115 700 117
rect 702 115 704 117
rect 698 113 704 115
rect 702 110 704 113
rect 722 118 728 120
rect 722 116 724 118
rect 726 116 728 118
rect 722 114 728 116
rect 732 118 738 120
rect 732 116 734 118
rect 736 116 738 118
rect 732 114 738 116
rect 722 111 724 114
rect 651 108 653 110
rect 655 108 657 110
rect 651 106 657 108
rect 637 103 639 106
rect 617 88 619 92
rect 627 85 629 90
rect 637 85 639 90
rect 597 79 599 83
rect 682 88 684 92
rect 692 88 694 92
rect 666 79 668 83
rect 735 104 737 114
rect 742 113 744 123
rect 762 120 764 125
rect 775 120 777 125
rect 762 118 768 120
rect 762 116 764 118
rect 766 116 768 118
rect 762 114 768 116
rect 772 118 778 120
rect 772 116 774 118
rect 776 116 778 118
rect 772 114 778 116
rect 742 111 748 113
rect 742 109 744 111
rect 746 109 748 111
rect 762 110 764 114
rect 742 107 748 109
rect 742 104 744 107
rect 722 88 724 93
rect 702 79 704 83
rect 772 103 774 114
rect 782 112 784 125
rect 867 134 869 138
rect 880 136 882 141
rect 887 136 889 141
rect 911 145 936 147
rect 911 137 913 145
rect 924 137 926 141
rect 934 137 936 145
rect 944 140 946 145
rect 951 140 953 145
rect 819 125 821 128
rect 812 123 821 125
rect 829 124 831 128
rect 839 125 841 128
rect 803 115 805 123
rect 812 121 814 123
rect 816 121 821 123
rect 812 119 821 121
rect 837 123 841 125
rect 837 120 839 123
rect 819 115 821 119
rect 833 118 839 120
rect 846 119 848 128
rect 908 135 913 137
rect 908 132 910 135
rect 867 120 869 125
rect 880 120 882 125
rect 833 116 835 118
rect 837 116 839 118
rect 800 113 813 115
rect 819 113 829 115
rect 833 114 839 116
rect 800 112 802 113
rect 782 110 788 112
rect 782 108 784 110
rect 786 108 788 110
rect 782 106 788 108
rect 796 110 802 112
rect 811 110 813 113
rect 827 110 829 113
rect 837 110 839 114
rect 843 117 849 119
rect 843 115 845 117
rect 847 115 849 117
rect 843 113 849 115
rect 847 110 849 113
rect 867 118 873 120
rect 867 116 869 118
rect 871 116 873 118
rect 867 114 873 116
rect 877 118 883 120
rect 877 116 879 118
rect 881 116 883 118
rect 877 114 883 116
rect 867 110 869 114
rect 796 108 798 110
rect 800 108 802 110
rect 796 106 802 108
rect 782 103 784 106
rect 762 88 764 92
rect 772 85 774 90
rect 782 85 784 90
rect 735 79 737 83
rect 742 79 744 83
rect 827 88 829 92
rect 837 88 839 92
rect 811 79 813 83
rect 877 103 879 114
rect 887 112 889 125
rect 972 132 974 137
rect 924 125 926 128
rect 917 123 926 125
rect 934 124 936 128
rect 944 125 946 128
rect 908 115 910 123
rect 917 121 919 123
rect 921 121 926 123
rect 917 119 926 121
rect 942 123 946 125
rect 942 120 944 123
rect 924 115 926 119
rect 938 118 944 120
rect 951 119 953 128
rect 982 129 984 134
rect 992 129 994 134
rect 1012 134 1014 138
rect 1025 136 1027 141
rect 1032 136 1034 141
rect 1056 145 1081 147
rect 1056 137 1058 145
rect 1069 137 1071 141
rect 1079 137 1081 145
rect 1089 140 1091 145
rect 1096 140 1098 145
rect 1053 135 1058 137
rect 1053 132 1055 135
rect 972 120 974 123
rect 982 120 984 123
rect 938 116 940 118
rect 942 116 944 118
rect 905 113 918 115
rect 924 113 934 115
rect 938 114 944 116
rect 905 112 907 113
rect 887 110 893 112
rect 887 108 889 110
rect 891 108 893 110
rect 887 106 893 108
rect 901 110 907 112
rect 916 110 918 113
rect 932 110 934 113
rect 942 110 944 114
rect 948 117 954 119
rect 948 115 950 117
rect 952 115 954 117
rect 948 113 954 115
rect 952 110 954 113
rect 972 118 978 120
rect 972 116 974 118
rect 976 116 978 118
rect 972 114 978 116
rect 982 118 988 120
rect 982 116 984 118
rect 986 116 988 118
rect 982 114 988 116
rect 972 111 974 114
rect 901 108 903 110
rect 905 108 907 110
rect 901 106 907 108
rect 887 103 889 106
rect 867 88 869 92
rect 877 85 879 90
rect 887 85 889 90
rect 847 79 849 83
rect 932 88 934 92
rect 942 88 944 92
rect 916 79 918 83
rect 985 104 987 114
rect 992 113 994 123
rect 1012 120 1014 125
rect 1025 120 1027 125
rect 1012 118 1018 120
rect 1012 116 1014 118
rect 1016 116 1018 118
rect 1012 114 1018 116
rect 1022 118 1028 120
rect 1022 116 1024 118
rect 1026 116 1028 118
rect 1022 114 1028 116
rect 992 111 998 113
rect 992 109 994 111
rect 996 109 998 111
rect 1012 110 1014 114
rect 992 107 998 109
rect 992 104 994 107
rect 972 88 974 93
rect 952 79 954 83
rect 1022 103 1024 114
rect 1032 112 1034 125
rect 1117 134 1119 138
rect 1130 136 1132 141
rect 1137 136 1139 141
rect 1161 145 1186 147
rect 1161 137 1163 145
rect 1174 137 1176 141
rect 1184 137 1186 145
rect 1194 140 1196 145
rect 1201 140 1203 145
rect 1069 125 1071 128
rect 1062 123 1071 125
rect 1079 124 1081 128
rect 1089 125 1091 128
rect 1053 115 1055 123
rect 1062 121 1064 123
rect 1066 121 1071 123
rect 1062 119 1071 121
rect 1087 123 1091 125
rect 1087 120 1089 123
rect 1069 115 1071 119
rect 1083 118 1089 120
rect 1096 119 1098 128
rect 1158 135 1163 137
rect 1158 132 1160 135
rect 1117 120 1119 125
rect 1130 120 1132 125
rect 1083 116 1085 118
rect 1087 116 1089 118
rect 1050 113 1063 115
rect 1069 113 1079 115
rect 1083 114 1089 116
rect 1050 112 1052 113
rect 1032 110 1038 112
rect 1032 108 1034 110
rect 1036 108 1038 110
rect 1032 106 1038 108
rect 1046 110 1052 112
rect 1061 110 1063 113
rect 1077 110 1079 113
rect 1087 110 1089 114
rect 1093 117 1099 119
rect 1093 115 1095 117
rect 1097 115 1099 117
rect 1093 113 1099 115
rect 1097 110 1099 113
rect 1117 118 1123 120
rect 1117 116 1119 118
rect 1121 116 1123 118
rect 1117 114 1123 116
rect 1127 118 1133 120
rect 1127 116 1129 118
rect 1131 116 1133 118
rect 1127 114 1133 116
rect 1117 110 1119 114
rect 1046 108 1048 110
rect 1050 108 1052 110
rect 1046 106 1052 108
rect 1032 103 1034 106
rect 1012 88 1014 92
rect 1022 85 1024 90
rect 1032 85 1034 90
rect 985 79 987 83
rect 992 79 994 83
rect 1077 88 1079 92
rect 1087 88 1089 92
rect 1061 79 1063 83
rect 1127 103 1129 114
rect 1137 112 1139 125
rect 1174 125 1176 128
rect 1167 123 1176 125
rect 1184 124 1186 128
rect 1194 125 1196 128
rect 1158 115 1160 123
rect 1167 121 1169 123
rect 1171 121 1176 123
rect 1167 119 1176 121
rect 1192 123 1196 125
rect 1192 120 1194 123
rect 1174 115 1176 119
rect 1188 118 1194 120
rect 1201 119 1203 128
rect 1188 116 1190 118
rect 1192 116 1194 118
rect 1155 113 1168 115
rect 1174 113 1184 115
rect 1188 114 1194 116
rect 1155 112 1157 113
rect 1137 110 1143 112
rect 1137 108 1139 110
rect 1141 108 1143 110
rect 1137 106 1143 108
rect 1151 110 1157 112
rect 1166 110 1168 113
rect 1182 110 1184 113
rect 1192 110 1194 114
rect 1198 117 1204 119
rect 1198 115 1200 117
rect 1202 115 1204 117
rect 1198 113 1204 115
rect 1202 110 1204 113
rect 1151 108 1153 110
rect 1155 108 1157 110
rect 1151 106 1157 108
rect 1137 103 1139 106
rect 1117 88 1119 92
rect 1127 85 1129 90
rect 1137 85 1139 90
rect 1097 79 1099 83
rect 1182 88 1184 92
rect 1192 88 1194 92
rect 1166 79 1168 83
rect 1202 79 1204 83
rect 27 71 29 75
rect 34 71 36 75
rect 14 61 16 66
rect 103 71 105 75
rect 54 62 56 66
rect 64 64 66 69
rect 74 64 76 69
rect 14 40 16 43
rect 27 40 29 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 31 16 34
rect 24 31 26 34
rect 34 31 36 41
rect 54 40 56 44
rect 64 40 66 51
rect 74 48 76 51
rect 74 46 80 48
rect 74 44 76 46
rect 78 44 80 46
rect 74 42 80 44
rect 88 46 94 48
rect 88 44 90 46
rect 92 44 94 46
rect 139 71 141 75
rect 119 62 121 66
rect 129 62 131 66
rect 208 71 210 75
rect 159 62 161 66
rect 169 64 171 69
rect 179 64 181 69
rect 88 42 94 44
rect 54 38 60 40
rect 54 36 56 38
rect 58 36 60 38
rect 54 34 60 36
rect 64 38 70 40
rect 64 36 66 38
rect 68 36 70 38
rect 64 34 70 36
rect 54 29 56 34
rect 67 29 69 34
rect 74 29 76 42
rect 92 41 94 42
rect 103 41 105 44
rect 119 41 121 44
rect 92 39 105 41
rect 111 39 121 41
rect 129 40 131 44
rect 139 41 141 44
rect 95 31 97 39
rect 111 35 113 39
rect 104 33 113 35
rect 125 38 131 40
rect 125 36 127 38
rect 129 36 131 38
rect 125 34 131 36
rect 135 39 141 41
rect 135 37 137 39
rect 139 37 141 39
rect 135 35 141 37
rect 159 40 161 44
rect 169 40 171 51
rect 179 48 181 51
rect 179 46 185 48
rect 179 44 181 46
rect 183 44 185 46
rect 179 42 185 44
rect 193 46 199 48
rect 193 44 195 46
rect 197 44 199 46
rect 244 71 246 75
rect 224 62 226 66
rect 234 62 236 66
rect 277 71 279 75
rect 284 71 286 75
rect 264 61 266 66
rect 193 42 199 44
rect 159 38 165 40
rect 159 36 161 38
rect 163 36 165 38
rect 104 31 106 33
rect 108 31 113 33
rect 14 17 16 22
rect 24 20 26 25
rect 34 20 36 25
rect 54 16 56 20
rect 104 29 113 31
rect 129 31 131 34
rect 111 26 113 29
rect 121 26 123 30
rect 129 29 133 31
rect 131 26 133 29
rect 138 26 140 35
rect 159 34 165 36
rect 169 38 175 40
rect 169 36 171 38
rect 173 36 175 38
rect 169 34 175 36
rect 159 29 161 34
rect 172 29 174 34
rect 179 29 181 42
rect 197 41 199 42
rect 208 41 210 44
rect 224 41 226 44
rect 197 39 210 41
rect 216 39 226 41
rect 234 40 236 44
rect 244 41 246 44
rect 353 71 355 75
rect 304 62 306 66
rect 314 64 316 69
rect 324 64 326 69
rect 200 31 202 39
rect 216 35 218 39
rect 209 33 218 35
rect 230 38 236 40
rect 230 36 232 38
rect 234 36 236 38
rect 230 34 236 36
rect 240 39 246 41
rect 240 37 242 39
rect 244 37 246 39
rect 240 35 246 37
rect 264 40 266 43
rect 277 40 279 50
rect 284 47 286 50
rect 284 45 290 47
rect 284 43 286 45
rect 288 43 290 45
rect 284 41 290 43
rect 264 38 270 40
rect 264 36 266 38
rect 268 36 270 38
rect 209 31 211 33
rect 213 31 218 33
rect 95 19 97 22
rect 67 13 69 18
rect 74 13 76 18
rect 95 17 100 19
rect 98 9 100 17
rect 111 13 113 17
rect 121 9 123 17
rect 159 16 161 20
rect 209 29 218 31
rect 234 31 236 34
rect 216 26 218 29
rect 226 26 228 30
rect 234 29 238 31
rect 236 26 238 29
rect 243 26 245 35
rect 264 34 270 36
rect 274 38 280 40
rect 274 36 276 38
rect 278 36 280 38
rect 274 34 280 36
rect 264 31 266 34
rect 274 31 276 34
rect 284 31 286 41
rect 304 40 306 44
rect 314 40 316 51
rect 324 48 326 51
rect 324 46 330 48
rect 324 44 326 46
rect 328 44 330 46
rect 324 42 330 44
rect 338 46 344 48
rect 338 44 340 46
rect 342 44 344 46
rect 389 71 391 75
rect 369 62 371 66
rect 379 62 381 66
rect 458 71 460 75
rect 409 62 411 66
rect 419 64 421 69
rect 429 64 431 69
rect 338 42 344 44
rect 304 38 310 40
rect 304 36 306 38
rect 308 36 310 38
rect 304 34 310 36
rect 314 38 320 40
rect 314 36 316 38
rect 318 36 320 38
rect 314 34 320 36
rect 200 19 202 22
rect 131 9 133 14
rect 138 9 140 14
rect 98 7 123 9
rect 172 13 174 18
rect 179 13 181 18
rect 200 17 205 19
rect 203 9 205 17
rect 216 13 218 17
rect 226 9 228 17
rect 304 29 306 34
rect 317 29 319 34
rect 324 29 326 42
rect 342 41 344 42
rect 353 41 355 44
rect 369 41 371 44
rect 342 39 355 41
rect 361 39 371 41
rect 379 40 381 44
rect 389 41 391 44
rect 345 31 347 39
rect 361 35 363 39
rect 354 33 363 35
rect 375 38 381 40
rect 375 36 377 38
rect 379 36 381 38
rect 375 34 381 36
rect 385 39 391 41
rect 385 37 387 39
rect 389 37 391 39
rect 385 35 391 37
rect 409 40 411 44
rect 419 40 421 51
rect 429 48 431 51
rect 429 46 435 48
rect 429 44 431 46
rect 433 44 435 46
rect 429 42 435 44
rect 443 46 449 48
rect 443 44 445 46
rect 447 44 449 46
rect 494 71 496 75
rect 474 62 476 66
rect 484 62 486 66
rect 527 71 529 75
rect 534 71 536 75
rect 514 61 516 66
rect 443 42 449 44
rect 409 38 415 40
rect 409 36 411 38
rect 413 36 415 38
rect 354 31 356 33
rect 358 31 363 33
rect 264 17 266 22
rect 274 20 276 25
rect 284 20 286 25
rect 236 9 238 14
rect 243 9 245 14
rect 203 7 228 9
rect 304 16 306 20
rect 354 29 363 31
rect 379 31 381 34
rect 361 26 363 29
rect 371 26 373 30
rect 379 29 383 31
rect 381 26 383 29
rect 388 26 390 35
rect 409 34 415 36
rect 419 38 425 40
rect 419 36 421 38
rect 423 36 425 38
rect 419 34 425 36
rect 409 29 411 34
rect 422 29 424 34
rect 429 29 431 42
rect 447 41 449 42
rect 458 41 460 44
rect 474 41 476 44
rect 447 39 460 41
rect 466 39 476 41
rect 484 40 486 44
rect 494 41 496 44
rect 603 71 605 75
rect 554 62 556 66
rect 564 64 566 69
rect 574 64 576 69
rect 450 31 452 39
rect 466 35 468 39
rect 459 33 468 35
rect 480 38 486 40
rect 480 36 482 38
rect 484 36 486 38
rect 480 34 486 36
rect 490 39 496 41
rect 490 37 492 39
rect 494 37 496 39
rect 490 35 496 37
rect 514 40 516 43
rect 527 40 529 50
rect 534 47 536 50
rect 534 45 540 47
rect 534 43 536 45
rect 538 43 540 45
rect 534 41 540 43
rect 514 38 520 40
rect 514 36 516 38
rect 518 36 520 38
rect 459 31 461 33
rect 463 31 468 33
rect 345 19 347 22
rect 317 13 319 18
rect 324 13 326 18
rect 345 17 350 19
rect 348 9 350 17
rect 361 13 363 17
rect 371 9 373 17
rect 409 16 411 20
rect 459 29 468 31
rect 484 31 486 34
rect 466 26 468 29
rect 476 26 478 30
rect 484 29 488 31
rect 486 26 488 29
rect 493 26 495 35
rect 514 34 520 36
rect 524 38 530 40
rect 524 36 526 38
rect 528 36 530 38
rect 524 34 530 36
rect 514 31 516 34
rect 524 31 526 34
rect 534 31 536 41
rect 554 40 556 44
rect 564 40 566 51
rect 574 48 576 51
rect 574 46 580 48
rect 574 44 576 46
rect 578 44 580 46
rect 574 42 580 44
rect 588 46 594 48
rect 588 44 590 46
rect 592 44 594 46
rect 639 71 641 75
rect 619 62 621 66
rect 629 62 631 66
rect 708 71 710 75
rect 659 62 661 66
rect 669 64 671 69
rect 679 64 681 69
rect 588 42 594 44
rect 554 38 560 40
rect 554 36 556 38
rect 558 36 560 38
rect 554 34 560 36
rect 564 38 570 40
rect 564 36 566 38
rect 568 36 570 38
rect 564 34 570 36
rect 450 19 452 22
rect 381 9 383 14
rect 388 9 390 14
rect 348 7 373 9
rect 422 13 424 18
rect 429 13 431 18
rect 450 17 455 19
rect 453 9 455 17
rect 466 13 468 17
rect 476 9 478 17
rect 554 29 556 34
rect 567 29 569 34
rect 574 29 576 42
rect 592 41 594 42
rect 603 41 605 44
rect 619 41 621 44
rect 592 39 605 41
rect 611 39 621 41
rect 629 40 631 44
rect 639 41 641 44
rect 595 31 597 39
rect 611 35 613 39
rect 604 33 613 35
rect 625 38 631 40
rect 625 36 627 38
rect 629 36 631 38
rect 625 34 631 36
rect 635 39 641 41
rect 635 37 637 39
rect 639 37 641 39
rect 635 35 641 37
rect 659 40 661 44
rect 669 40 671 51
rect 679 48 681 51
rect 679 46 685 48
rect 679 44 681 46
rect 683 44 685 46
rect 679 42 685 44
rect 693 46 699 48
rect 693 44 695 46
rect 697 44 699 46
rect 744 71 746 75
rect 724 62 726 66
rect 734 62 736 66
rect 777 71 779 75
rect 784 71 786 75
rect 764 61 766 66
rect 693 42 699 44
rect 659 38 665 40
rect 659 36 661 38
rect 663 36 665 38
rect 604 31 606 33
rect 608 31 613 33
rect 514 17 516 22
rect 524 20 526 25
rect 534 20 536 25
rect 486 9 488 14
rect 493 9 495 14
rect 453 7 478 9
rect 554 16 556 20
rect 604 29 613 31
rect 629 31 631 34
rect 611 26 613 29
rect 621 26 623 30
rect 629 29 633 31
rect 631 26 633 29
rect 638 26 640 35
rect 659 34 665 36
rect 669 38 675 40
rect 669 36 671 38
rect 673 36 675 38
rect 669 34 675 36
rect 659 29 661 34
rect 672 29 674 34
rect 679 29 681 42
rect 697 41 699 42
rect 708 41 710 44
rect 724 41 726 44
rect 697 39 710 41
rect 716 39 726 41
rect 734 40 736 44
rect 744 41 746 44
rect 853 71 855 75
rect 804 62 806 66
rect 814 64 816 69
rect 824 64 826 69
rect 700 31 702 39
rect 716 35 718 39
rect 709 33 718 35
rect 730 38 736 40
rect 730 36 732 38
rect 734 36 736 38
rect 730 34 736 36
rect 740 39 746 41
rect 740 37 742 39
rect 744 37 746 39
rect 740 35 746 37
rect 764 40 766 43
rect 777 40 779 50
rect 784 47 786 50
rect 784 45 790 47
rect 784 43 786 45
rect 788 43 790 45
rect 784 41 790 43
rect 764 38 770 40
rect 764 36 766 38
rect 768 36 770 38
rect 709 31 711 33
rect 713 31 718 33
rect 595 19 597 22
rect 567 13 569 18
rect 574 13 576 18
rect 595 17 600 19
rect 598 9 600 17
rect 611 13 613 17
rect 621 9 623 17
rect 659 16 661 20
rect 709 29 718 31
rect 734 31 736 34
rect 716 26 718 29
rect 726 26 728 30
rect 734 29 738 31
rect 736 26 738 29
rect 743 26 745 35
rect 764 34 770 36
rect 774 38 780 40
rect 774 36 776 38
rect 778 36 780 38
rect 774 34 780 36
rect 764 31 766 34
rect 774 31 776 34
rect 784 31 786 41
rect 804 40 806 44
rect 814 40 816 51
rect 824 48 826 51
rect 824 46 830 48
rect 824 44 826 46
rect 828 44 830 46
rect 824 42 830 44
rect 838 46 844 48
rect 838 44 840 46
rect 842 44 844 46
rect 889 71 891 75
rect 869 62 871 66
rect 879 62 881 66
rect 958 71 960 75
rect 909 62 911 66
rect 919 64 921 69
rect 929 64 931 69
rect 838 42 844 44
rect 804 38 810 40
rect 804 36 806 38
rect 808 36 810 38
rect 804 34 810 36
rect 814 38 820 40
rect 814 36 816 38
rect 818 36 820 38
rect 814 34 820 36
rect 700 19 702 22
rect 631 9 633 14
rect 638 9 640 14
rect 598 7 623 9
rect 672 13 674 18
rect 679 13 681 18
rect 700 17 705 19
rect 703 9 705 17
rect 716 13 718 17
rect 726 9 728 17
rect 804 29 806 34
rect 817 29 819 34
rect 824 29 826 42
rect 842 41 844 42
rect 853 41 855 44
rect 869 41 871 44
rect 842 39 855 41
rect 861 39 871 41
rect 879 40 881 44
rect 889 41 891 44
rect 845 31 847 39
rect 861 35 863 39
rect 854 33 863 35
rect 875 38 881 40
rect 875 36 877 38
rect 879 36 881 38
rect 875 34 881 36
rect 885 39 891 41
rect 885 37 887 39
rect 889 37 891 39
rect 885 35 891 37
rect 909 40 911 44
rect 919 40 921 51
rect 929 48 931 51
rect 929 46 935 48
rect 929 44 931 46
rect 933 44 935 46
rect 929 42 935 44
rect 943 46 949 48
rect 943 44 945 46
rect 947 44 949 46
rect 994 71 996 75
rect 974 62 976 66
rect 984 62 986 66
rect 943 42 949 44
rect 909 38 915 40
rect 909 36 911 38
rect 913 36 915 38
rect 854 31 856 33
rect 858 31 863 33
rect 764 17 766 22
rect 774 20 776 25
rect 784 20 786 25
rect 736 9 738 14
rect 743 9 745 14
rect 703 7 728 9
rect 804 16 806 20
rect 854 29 863 31
rect 879 31 881 34
rect 861 26 863 29
rect 871 26 873 30
rect 879 29 883 31
rect 881 26 883 29
rect 888 26 890 35
rect 909 34 915 36
rect 919 38 925 40
rect 919 36 921 38
rect 923 36 925 38
rect 919 34 925 36
rect 909 29 911 34
rect 922 29 924 34
rect 929 29 931 42
rect 947 41 949 42
rect 958 41 960 44
rect 974 41 976 44
rect 947 39 960 41
rect 966 39 976 41
rect 984 40 986 44
rect 994 41 996 44
rect 950 31 952 39
rect 966 35 968 39
rect 959 33 968 35
rect 980 38 986 40
rect 980 36 982 38
rect 984 36 986 38
rect 980 34 986 36
rect 990 39 996 41
rect 990 37 992 39
rect 994 37 996 39
rect 990 35 996 37
rect 959 31 961 33
rect 963 31 968 33
rect 845 19 847 22
rect 817 13 819 18
rect 824 13 826 18
rect 845 17 850 19
rect 848 9 850 17
rect 861 13 863 17
rect 871 9 873 17
rect 909 16 911 20
rect 959 29 968 31
rect 984 31 986 34
rect 966 26 968 29
rect 976 26 978 30
rect 984 29 988 31
rect 986 26 988 29
rect 993 26 995 35
rect 950 19 952 22
rect 881 9 883 14
rect 888 9 890 14
rect 848 7 873 9
rect 922 13 924 18
rect 929 13 931 18
rect 950 17 955 19
rect 953 9 955 17
rect 966 13 968 17
rect 976 9 978 17
rect 986 9 988 14
rect 993 9 995 14
rect 953 7 978 9
<< ndif >>
rect 32 413 39 415
rect 32 411 35 413
rect 37 411 39 413
rect 32 405 39 411
rect 72 413 79 415
rect 72 411 75 413
rect 77 411 79 413
rect 14 403 21 405
rect 14 401 16 403
rect 18 401 21 403
rect 14 399 21 401
rect 16 394 21 399
rect 23 394 28 405
rect 30 403 39 405
rect 72 405 79 411
rect 101 413 107 415
rect 514 415 521 417
rect 101 411 103 413
rect 105 411 107 413
rect 101 409 107 411
rect 54 403 61 405
rect 30 394 41 403
rect 43 401 50 403
rect 43 399 46 401
rect 48 399 50 401
rect 54 401 56 403
rect 58 401 61 403
rect 54 399 61 401
rect 43 397 50 399
rect 43 394 48 397
rect 56 394 61 399
rect 63 394 68 405
rect 70 403 79 405
rect 70 394 81 403
rect 83 401 90 403
rect 83 399 86 401
rect 88 399 90 401
rect 83 397 90 399
rect 101 397 109 409
rect 111 397 116 409
rect 118 406 123 409
rect 184 413 191 415
rect 184 411 187 413
rect 189 411 191 413
rect 118 403 126 406
rect 118 401 121 403
rect 123 401 126 403
rect 118 397 126 401
rect 128 401 136 406
rect 128 399 131 401
rect 133 399 136 401
rect 128 397 136 399
rect 138 404 147 406
rect 184 405 191 411
rect 514 413 517 415
rect 519 413 521 415
rect 514 407 521 413
rect 554 415 561 417
rect 554 413 557 415
rect 559 413 561 415
rect 138 402 143 404
rect 145 402 147 404
rect 138 401 147 402
rect 166 403 173 405
rect 166 401 168 403
rect 170 401 173 403
rect 138 397 152 401
rect 83 394 88 397
rect 147 392 152 397
rect 154 398 159 401
rect 166 399 173 401
rect 154 396 161 398
rect 154 394 157 396
rect 159 394 161 396
rect 168 394 173 399
rect 175 394 180 405
rect 182 403 191 405
rect 496 405 503 407
rect 496 403 498 405
rect 500 403 503 405
rect 182 394 193 403
rect 195 401 202 403
rect 496 401 503 403
rect 195 399 198 401
rect 200 399 202 401
rect 195 397 202 399
rect 195 394 200 397
rect 498 396 503 401
rect 505 396 510 407
rect 512 405 521 407
rect 554 407 561 413
rect 583 415 589 417
rect 583 413 585 415
rect 587 413 589 415
rect 583 411 589 413
rect 536 405 543 407
rect 512 396 523 405
rect 525 403 532 405
rect 525 401 528 403
rect 530 401 532 403
rect 536 403 538 405
rect 540 403 543 405
rect 536 401 543 403
rect 525 399 532 401
rect 525 396 530 399
rect 538 396 543 401
rect 545 396 550 407
rect 552 405 561 407
rect 552 396 563 405
rect 565 403 572 405
rect 565 401 568 403
rect 570 401 572 403
rect 565 399 572 401
rect 583 399 591 411
rect 593 399 598 411
rect 600 408 605 411
rect 666 415 673 417
rect 666 413 669 415
rect 671 413 673 415
rect 600 405 608 408
rect 600 403 603 405
rect 605 403 608 405
rect 600 399 608 403
rect 610 403 618 408
rect 610 401 613 403
rect 615 401 618 403
rect 610 399 618 401
rect 620 406 629 408
rect 666 407 673 413
rect 719 415 726 417
rect 719 413 722 415
rect 724 413 726 415
rect 620 404 625 406
rect 627 404 629 406
rect 620 403 629 404
rect 648 405 655 407
rect 648 403 650 405
rect 652 403 655 405
rect 620 399 634 403
rect 565 396 570 399
rect 154 392 161 394
rect 629 394 634 399
rect 636 400 641 403
rect 648 401 655 403
rect 636 398 643 400
rect 636 396 639 398
rect 641 396 643 398
rect 650 396 655 401
rect 657 396 662 407
rect 664 405 673 407
rect 719 407 726 413
rect 759 415 766 417
rect 759 413 762 415
rect 764 413 766 415
rect 701 405 708 407
rect 664 396 675 405
rect 677 403 684 405
rect 677 401 680 403
rect 682 401 684 403
rect 701 403 703 405
rect 705 403 708 405
rect 701 401 708 403
rect 677 399 684 401
rect 677 396 682 399
rect 703 396 708 401
rect 710 396 715 407
rect 717 405 726 407
rect 759 407 766 413
rect 788 415 794 417
rect 788 413 790 415
rect 792 413 794 415
rect 788 411 794 413
rect 741 405 748 407
rect 717 396 728 405
rect 730 403 737 405
rect 730 401 733 403
rect 735 401 737 403
rect 741 403 743 405
rect 745 403 748 405
rect 741 401 748 403
rect 730 399 737 401
rect 730 396 735 399
rect 743 396 748 401
rect 750 396 755 407
rect 757 405 766 407
rect 757 396 768 405
rect 770 403 777 405
rect 770 401 773 403
rect 775 401 777 403
rect 770 399 777 401
rect 788 399 796 411
rect 798 399 803 411
rect 805 408 810 411
rect 871 415 878 417
rect 871 413 874 415
rect 876 413 878 415
rect 805 405 813 408
rect 805 403 808 405
rect 810 403 813 405
rect 805 399 813 403
rect 815 403 823 408
rect 815 401 818 403
rect 820 401 823 403
rect 815 399 823 401
rect 825 406 834 408
rect 871 407 878 413
rect 825 404 830 406
rect 832 404 834 406
rect 825 403 834 404
rect 853 405 860 407
rect 853 403 855 405
rect 857 403 860 405
rect 825 399 839 403
rect 770 396 775 399
rect 636 394 643 396
rect 834 394 839 399
rect 841 400 846 403
rect 853 401 860 403
rect 841 398 848 400
rect 841 396 844 398
rect 846 396 848 398
rect 855 396 860 401
rect 862 396 867 407
rect 869 405 878 407
rect 869 396 880 405
rect 882 403 889 405
rect 882 401 885 403
rect 887 401 889 403
rect 882 399 889 401
rect 882 396 887 399
rect 841 394 848 396
rect 135 298 142 300
rect 16 295 21 298
rect 14 293 21 295
rect 14 291 16 293
rect 18 291 21 293
rect 14 289 21 291
rect 23 289 34 298
rect 25 287 34 289
rect 36 287 41 298
rect 43 293 48 298
rect 56 293 61 298
rect 43 291 50 293
rect 43 289 46 291
rect 48 289 50 291
rect 43 287 50 289
rect 54 291 61 293
rect 54 289 56 291
rect 58 289 61 291
rect 54 287 61 289
rect 63 287 68 298
rect 70 289 81 298
rect 83 295 88 298
rect 96 295 101 298
rect 83 293 90 295
rect 83 291 86 293
rect 88 291 90 293
rect 83 289 90 291
rect 94 293 101 295
rect 94 291 96 293
rect 98 291 101 293
rect 94 289 101 291
rect 103 289 114 298
rect 70 287 79 289
rect 25 281 32 287
rect 25 279 27 281
rect 29 279 32 281
rect 25 277 32 279
rect 72 281 79 287
rect 105 287 114 289
rect 116 287 121 298
rect 123 293 128 298
rect 135 296 137 298
rect 139 296 142 298
rect 135 294 142 296
rect 123 291 130 293
rect 137 291 142 294
rect 144 295 149 300
rect 617 300 624 302
rect 498 297 503 300
rect 496 295 503 297
rect 144 291 158 295
rect 123 289 126 291
rect 128 289 130 291
rect 123 287 130 289
rect 149 290 158 291
rect 149 288 151 290
rect 153 288 158 290
rect 72 279 75 281
rect 77 279 79 281
rect 72 277 79 279
rect 105 281 112 287
rect 149 286 158 288
rect 160 293 168 295
rect 160 291 163 293
rect 165 291 168 293
rect 160 286 168 291
rect 170 291 178 295
rect 170 289 173 291
rect 175 289 178 291
rect 170 286 178 289
rect 105 279 107 281
rect 109 279 112 281
rect 105 277 112 279
rect 173 283 178 286
rect 180 283 185 295
rect 187 283 195 295
rect 496 293 498 295
rect 500 293 503 295
rect 496 291 503 293
rect 505 291 516 300
rect 507 289 516 291
rect 518 289 523 300
rect 525 295 530 300
rect 538 295 543 300
rect 525 293 532 295
rect 525 291 528 293
rect 530 291 532 293
rect 525 289 532 291
rect 536 293 543 295
rect 536 291 538 293
rect 540 291 543 293
rect 536 289 543 291
rect 545 289 550 300
rect 552 291 563 300
rect 565 297 570 300
rect 578 297 583 300
rect 565 295 572 297
rect 565 293 568 295
rect 570 293 572 295
rect 565 291 572 293
rect 576 295 583 297
rect 576 293 578 295
rect 580 293 583 295
rect 576 291 583 293
rect 585 291 596 300
rect 552 289 561 291
rect 189 281 195 283
rect 189 279 191 281
rect 193 279 195 281
rect 507 283 514 289
rect 507 281 509 283
rect 511 281 514 283
rect 507 279 514 281
rect 554 283 561 289
rect 587 289 596 291
rect 598 289 603 300
rect 605 295 610 300
rect 617 298 619 300
rect 621 298 624 300
rect 617 296 624 298
rect 605 293 612 295
rect 619 293 624 296
rect 626 297 631 302
rect 822 300 829 302
rect 703 297 708 300
rect 626 293 640 297
rect 605 291 608 293
rect 610 291 612 293
rect 605 289 612 291
rect 631 292 640 293
rect 631 290 633 292
rect 635 290 640 292
rect 554 281 557 283
rect 559 281 561 283
rect 554 279 561 281
rect 587 283 594 289
rect 631 288 640 290
rect 642 295 650 297
rect 642 293 645 295
rect 647 293 650 295
rect 642 288 650 293
rect 652 293 660 297
rect 652 291 655 293
rect 657 291 660 293
rect 652 288 660 291
rect 587 281 589 283
rect 591 281 594 283
rect 587 279 594 281
rect 655 285 660 288
rect 662 285 667 297
rect 669 285 677 297
rect 701 295 708 297
rect 701 293 703 295
rect 705 293 708 295
rect 701 291 708 293
rect 710 291 721 300
rect 712 289 721 291
rect 723 289 728 300
rect 730 295 735 300
rect 743 295 748 300
rect 730 293 737 295
rect 730 291 733 293
rect 735 291 737 293
rect 730 289 737 291
rect 741 293 748 295
rect 741 291 743 293
rect 745 291 748 293
rect 741 289 748 291
rect 750 289 755 300
rect 757 291 768 300
rect 770 297 775 300
rect 783 297 788 300
rect 770 295 777 297
rect 770 293 773 295
rect 775 293 777 295
rect 770 291 777 293
rect 781 295 788 297
rect 781 293 783 295
rect 785 293 788 295
rect 781 291 788 293
rect 790 291 801 300
rect 757 289 766 291
rect 671 283 677 285
rect 671 281 673 283
rect 675 281 677 283
rect 189 277 195 279
rect 671 279 677 281
rect 712 283 719 289
rect 712 281 714 283
rect 716 281 719 283
rect 712 279 719 281
rect 759 283 766 289
rect 792 289 801 291
rect 803 289 808 300
rect 810 295 815 300
rect 822 298 824 300
rect 826 298 829 300
rect 822 296 829 298
rect 810 293 817 295
rect 824 293 829 296
rect 831 297 836 302
rect 1040 297 1047 299
rect 831 293 845 297
rect 810 291 813 293
rect 815 291 817 293
rect 810 289 817 291
rect 836 292 845 293
rect 836 290 838 292
rect 840 290 845 292
rect 759 281 762 283
rect 764 281 766 283
rect 759 279 766 281
rect 792 283 799 289
rect 836 288 845 290
rect 847 295 855 297
rect 847 293 850 295
rect 852 293 855 295
rect 847 288 855 293
rect 857 293 865 297
rect 857 291 860 293
rect 862 291 865 293
rect 857 288 865 291
rect 792 281 794 283
rect 796 281 799 283
rect 792 279 799 281
rect 860 285 865 288
rect 867 285 872 297
rect 874 285 882 297
rect 1040 295 1043 297
rect 1045 295 1047 297
rect 1040 289 1047 295
rect 1080 297 1087 299
rect 1080 295 1083 297
rect 1085 295 1087 297
rect 876 283 882 285
rect 1022 287 1029 289
rect 1022 285 1024 287
rect 1026 285 1029 287
rect 1022 283 1029 285
rect 876 281 878 283
rect 880 281 882 283
rect 876 279 882 281
rect 1024 278 1029 283
rect 1031 278 1036 289
rect 1038 287 1047 289
rect 1080 289 1087 295
rect 1109 297 1115 299
rect 1109 295 1111 297
rect 1113 295 1115 297
rect 1109 293 1115 295
rect 1062 287 1069 289
rect 1038 278 1049 287
rect 1051 285 1058 287
rect 1051 283 1054 285
rect 1056 283 1058 285
rect 1062 285 1064 287
rect 1066 285 1069 287
rect 1062 283 1069 285
rect 1051 281 1058 283
rect 1051 278 1056 281
rect 1064 278 1069 283
rect 1071 278 1076 289
rect 1078 287 1087 289
rect 1078 278 1089 287
rect 1091 285 1098 287
rect 1091 283 1094 285
rect 1096 283 1098 285
rect 1091 281 1098 283
rect 1109 281 1117 293
rect 1119 281 1124 293
rect 1126 290 1131 293
rect 1192 297 1199 299
rect 1192 295 1195 297
rect 1197 295 1199 297
rect 1126 287 1134 290
rect 1126 285 1129 287
rect 1131 285 1134 287
rect 1126 281 1134 285
rect 1136 285 1144 290
rect 1136 283 1139 285
rect 1141 283 1144 285
rect 1136 281 1144 283
rect 1146 288 1155 290
rect 1192 289 1199 295
rect 1146 286 1151 288
rect 1153 286 1155 288
rect 1146 285 1155 286
rect 1174 287 1181 289
rect 1174 285 1176 287
rect 1178 285 1181 287
rect 1146 281 1160 285
rect 1091 278 1096 281
rect 1155 276 1160 281
rect 1162 282 1167 285
rect 1174 283 1181 285
rect 1162 280 1169 282
rect 1162 278 1165 280
rect 1167 278 1169 280
rect 1176 278 1181 283
rect 1183 278 1188 289
rect 1190 287 1199 289
rect 1190 278 1201 287
rect 1203 285 1210 287
rect 1203 283 1206 285
rect 1208 283 1210 285
rect 1203 281 1210 283
rect 1203 278 1208 281
rect 1162 276 1169 278
rect 1 182 8 184
rect 1 180 3 182
rect 5 180 8 182
rect 1 178 8 180
rect 3 175 8 178
rect 10 178 18 184
rect 20 182 28 184
rect 20 180 23 182
rect 25 180 28 182
rect 20 178 28 180
rect 30 178 37 184
rect 82 182 89 184
rect 43 179 48 182
rect 10 175 16 178
rect 12 171 16 175
rect 32 171 37 178
rect 41 177 48 179
rect 41 175 43 177
rect 45 175 48 177
rect 41 173 48 175
rect 50 173 61 182
rect 12 169 18 171
rect 12 167 14 169
rect 16 167 18 169
rect 12 165 18 167
rect 31 169 37 171
rect 52 171 61 173
rect 63 171 68 182
rect 70 177 75 182
rect 82 180 84 182
rect 86 180 89 182
rect 82 178 89 180
rect 70 175 77 177
rect 84 175 89 178
rect 91 179 96 184
rect 187 182 194 184
rect 148 179 153 182
rect 91 175 105 179
rect 70 173 73 175
rect 75 173 77 175
rect 70 171 77 173
rect 96 174 105 175
rect 96 172 98 174
rect 100 172 105 174
rect 31 167 33 169
rect 35 167 37 169
rect 31 165 37 167
rect 52 165 59 171
rect 96 170 105 172
rect 107 177 115 179
rect 107 175 110 177
rect 112 175 115 177
rect 107 170 115 175
rect 117 175 125 179
rect 117 173 120 175
rect 122 173 125 175
rect 117 170 125 173
rect 52 163 54 165
rect 56 163 59 165
rect 52 161 59 163
rect 120 167 125 170
rect 127 167 132 179
rect 134 167 142 179
rect 146 177 153 179
rect 146 175 148 177
rect 150 175 153 177
rect 146 173 153 175
rect 155 173 166 182
rect 157 171 166 173
rect 168 171 173 182
rect 175 177 180 182
rect 187 180 189 182
rect 191 180 194 182
rect 187 178 194 180
rect 175 175 182 177
rect 189 175 194 178
rect 196 179 201 184
rect 251 182 258 184
rect 251 180 253 182
rect 255 180 258 182
rect 196 175 210 179
rect 175 173 178 175
rect 180 173 182 175
rect 175 171 182 173
rect 201 174 210 175
rect 201 172 203 174
rect 205 172 210 174
rect 136 165 142 167
rect 136 163 138 165
rect 140 163 142 165
rect 136 161 142 163
rect 157 165 164 171
rect 201 170 210 172
rect 212 177 220 179
rect 212 175 215 177
rect 217 175 220 177
rect 212 170 220 175
rect 222 175 230 179
rect 222 173 225 175
rect 227 173 230 175
rect 222 170 230 173
rect 157 163 159 165
rect 161 163 164 165
rect 157 161 164 163
rect 225 167 230 170
rect 232 167 237 179
rect 239 167 247 179
rect 251 178 258 180
rect 253 175 258 178
rect 260 178 268 184
rect 270 182 278 184
rect 270 180 273 182
rect 275 180 278 182
rect 270 178 278 180
rect 280 178 287 184
rect 332 182 339 184
rect 293 179 298 182
rect 260 175 266 178
rect 262 171 266 175
rect 282 171 287 178
rect 291 177 298 179
rect 291 175 293 177
rect 295 175 298 177
rect 291 173 298 175
rect 300 173 311 182
rect 262 169 268 171
rect 262 167 264 169
rect 266 167 268 169
rect 241 165 247 167
rect 241 163 243 165
rect 245 163 247 165
rect 241 161 247 163
rect 262 165 268 167
rect 281 169 287 171
rect 302 171 311 173
rect 313 171 318 182
rect 320 177 325 182
rect 332 180 334 182
rect 336 180 339 182
rect 332 178 339 180
rect 320 175 327 177
rect 334 175 339 178
rect 341 179 346 184
rect 437 182 444 184
rect 398 179 403 182
rect 341 175 355 179
rect 320 173 323 175
rect 325 173 327 175
rect 320 171 327 173
rect 346 174 355 175
rect 346 172 348 174
rect 350 172 355 174
rect 281 167 283 169
rect 285 167 287 169
rect 281 165 287 167
rect 302 165 309 171
rect 346 170 355 172
rect 357 177 365 179
rect 357 175 360 177
rect 362 175 365 177
rect 357 170 365 175
rect 367 175 375 179
rect 367 173 370 175
rect 372 173 375 175
rect 367 170 375 173
rect 302 163 304 165
rect 306 163 309 165
rect 302 161 309 163
rect 370 167 375 170
rect 377 167 382 179
rect 384 167 392 179
rect 396 177 403 179
rect 396 175 398 177
rect 400 175 403 177
rect 396 173 403 175
rect 405 173 416 182
rect 407 171 416 173
rect 418 171 423 182
rect 425 177 430 182
rect 437 180 439 182
rect 441 180 444 182
rect 437 178 444 180
rect 425 175 432 177
rect 439 175 444 178
rect 446 179 451 184
rect 501 182 508 184
rect 501 180 503 182
rect 505 180 508 182
rect 446 175 460 179
rect 425 173 428 175
rect 430 173 432 175
rect 425 171 432 173
rect 451 174 460 175
rect 451 172 453 174
rect 455 172 460 174
rect 386 165 392 167
rect 386 163 388 165
rect 390 163 392 165
rect 386 161 392 163
rect 407 165 414 171
rect 451 170 460 172
rect 462 177 470 179
rect 462 175 465 177
rect 467 175 470 177
rect 462 170 470 175
rect 472 175 480 179
rect 472 173 475 175
rect 477 173 480 175
rect 472 170 480 173
rect 407 163 409 165
rect 411 163 414 165
rect 407 161 414 163
rect 475 167 480 170
rect 482 167 487 179
rect 489 167 497 179
rect 501 178 508 180
rect 503 175 508 178
rect 510 178 518 184
rect 520 182 528 184
rect 520 180 523 182
rect 525 180 528 182
rect 520 178 528 180
rect 530 178 537 184
rect 582 182 589 184
rect 543 179 548 182
rect 510 175 516 178
rect 512 171 516 175
rect 532 171 537 178
rect 541 177 548 179
rect 541 175 543 177
rect 545 175 548 177
rect 541 173 548 175
rect 550 173 561 182
rect 512 169 518 171
rect 512 167 514 169
rect 516 167 518 169
rect 491 165 497 167
rect 491 163 493 165
rect 495 163 497 165
rect 491 161 497 163
rect 512 165 518 167
rect 531 169 537 171
rect 552 171 561 173
rect 563 171 568 182
rect 570 177 575 182
rect 582 180 584 182
rect 586 180 589 182
rect 582 178 589 180
rect 570 175 577 177
rect 584 175 589 178
rect 591 179 596 184
rect 687 182 694 184
rect 648 179 653 182
rect 591 175 605 179
rect 570 173 573 175
rect 575 173 577 175
rect 570 171 577 173
rect 596 174 605 175
rect 596 172 598 174
rect 600 172 605 174
rect 531 167 533 169
rect 535 167 537 169
rect 531 165 537 167
rect 552 165 559 171
rect 596 170 605 172
rect 607 177 615 179
rect 607 175 610 177
rect 612 175 615 177
rect 607 170 615 175
rect 617 175 625 179
rect 617 173 620 175
rect 622 173 625 175
rect 617 170 625 173
rect 552 163 554 165
rect 556 163 559 165
rect 552 161 559 163
rect 620 167 625 170
rect 627 167 632 179
rect 634 167 642 179
rect 646 177 653 179
rect 646 175 648 177
rect 650 175 653 177
rect 646 173 653 175
rect 655 173 666 182
rect 657 171 666 173
rect 668 171 673 182
rect 675 177 680 182
rect 687 180 689 182
rect 691 180 694 182
rect 687 178 694 180
rect 675 175 682 177
rect 689 175 694 178
rect 696 179 701 184
rect 751 182 758 184
rect 751 180 753 182
rect 755 180 758 182
rect 696 175 710 179
rect 675 173 678 175
rect 680 173 682 175
rect 675 171 682 173
rect 701 174 710 175
rect 701 172 703 174
rect 705 172 710 174
rect 636 165 642 167
rect 636 163 638 165
rect 640 163 642 165
rect 636 161 642 163
rect 657 165 664 171
rect 701 170 710 172
rect 712 177 720 179
rect 712 175 715 177
rect 717 175 720 177
rect 712 170 720 175
rect 722 175 730 179
rect 722 173 725 175
rect 727 173 730 175
rect 722 170 730 173
rect 657 163 659 165
rect 661 163 664 165
rect 657 161 664 163
rect 725 167 730 170
rect 732 167 737 179
rect 739 167 747 179
rect 751 178 758 180
rect 753 175 758 178
rect 760 178 768 184
rect 770 182 778 184
rect 770 180 773 182
rect 775 180 778 182
rect 770 178 778 180
rect 780 178 787 184
rect 832 182 839 184
rect 793 179 798 182
rect 760 175 766 178
rect 762 171 766 175
rect 782 171 787 178
rect 791 177 798 179
rect 791 175 793 177
rect 795 175 798 177
rect 791 173 798 175
rect 800 173 811 182
rect 762 169 768 171
rect 762 167 764 169
rect 766 167 768 169
rect 741 165 747 167
rect 741 163 743 165
rect 745 163 747 165
rect 741 161 747 163
rect 762 165 768 167
rect 781 169 787 171
rect 802 171 811 173
rect 813 171 818 182
rect 820 177 825 182
rect 832 180 834 182
rect 836 180 839 182
rect 832 178 839 180
rect 820 175 827 177
rect 834 175 839 178
rect 841 179 846 184
rect 937 182 944 184
rect 898 179 903 182
rect 841 175 855 179
rect 820 173 823 175
rect 825 173 827 175
rect 820 171 827 173
rect 846 174 855 175
rect 846 172 848 174
rect 850 172 855 174
rect 781 167 783 169
rect 785 167 787 169
rect 781 165 787 167
rect 802 165 809 171
rect 846 170 855 172
rect 857 177 865 179
rect 857 175 860 177
rect 862 175 865 177
rect 857 170 865 175
rect 867 175 875 179
rect 867 173 870 175
rect 872 173 875 175
rect 867 170 875 173
rect 802 163 804 165
rect 806 163 809 165
rect 802 161 809 163
rect 870 167 875 170
rect 877 167 882 179
rect 884 167 892 179
rect 896 177 903 179
rect 896 175 898 177
rect 900 175 903 177
rect 896 173 903 175
rect 905 173 916 182
rect 907 171 916 173
rect 918 171 923 182
rect 925 177 930 182
rect 937 180 939 182
rect 941 180 944 182
rect 937 178 944 180
rect 925 175 932 177
rect 939 175 944 178
rect 946 179 951 184
rect 1143 182 1150 184
rect 1024 179 1029 182
rect 946 175 960 179
rect 925 173 928 175
rect 930 173 932 175
rect 925 171 932 173
rect 951 174 960 175
rect 951 172 953 174
rect 955 172 960 174
rect 886 165 892 167
rect 886 163 888 165
rect 890 163 892 165
rect 886 161 892 163
rect 907 165 914 171
rect 951 170 960 172
rect 962 177 970 179
rect 962 175 965 177
rect 967 175 970 177
rect 962 170 970 175
rect 972 175 980 179
rect 972 173 975 175
rect 977 173 980 175
rect 972 170 980 173
rect 907 163 909 165
rect 911 163 914 165
rect 907 161 914 163
rect 975 167 980 170
rect 982 167 987 179
rect 989 167 997 179
rect 1022 177 1029 179
rect 1022 175 1024 177
rect 1026 175 1029 177
rect 1022 173 1029 175
rect 1031 173 1042 182
rect 1033 171 1042 173
rect 1044 171 1049 182
rect 1051 177 1056 182
rect 1064 177 1069 182
rect 1051 175 1058 177
rect 1051 173 1054 175
rect 1056 173 1058 175
rect 1051 171 1058 173
rect 1062 175 1069 177
rect 1062 173 1064 175
rect 1066 173 1069 175
rect 1062 171 1069 173
rect 1071 171 1076 182
rect 1078 173 1089 182
rect 1091 179 1096 182
rect 1104 179 1109 182
rect 1091 177 1098 179
rect 1091 175 1094 177
rect 1096 175 1098 177
rect 1091 173 1098 175
rect 1102 177 1109 179
rect 1102 175 1104 177
rect 1106 175 1109 177
rect 1102 173 1109 175
rect 1111 173 1122 182
rect 1078 171 1087 173
rect 991 165 997 167
rect 991 163 993 165
rect 995 163 997 165
rect 991 161 997 163
rect 1033 165 1040 171
rect 1033 163 1035 165
rect 1037 163 1040 165
rect 1033 161 1040 163
rect 1080 165 1087 171
rect 1113 171 1122 173
rect 1124 171 1129 182
rect 1131 177 1136 182
rect 1143 180 1145 182
rect 1147 180 1150 182
rect 1143 178 1150 180
rect 1131 175 1138 177
rect 1145 175 1150 178
rect 1152 179 1157 184
rect 1152 175 1166 179
rect 1131 173 1134 175
rect 1136 173 1138 175
rect 1131 171 1138 173
rect 1157 174 1166 175
rect 1157 172 1159 174
rect 1161 172 1166 174
rect 1080 163 1083 165
rect 1085 163 1087 165
rect 1080 161 1087 163
rect 1113 165 1120 171
rect 1157 170 1166 172
rect 1168 177 1176 179
rect 1168 175 1171 177
rect 1173 175 1176 177
rect 1168 170 1176 175
rect 1178 175 1186 179
rect 1178 173 1181 175
rect 1183 173 1186 175
rect 1178 170 1186 173
rect 1113 163 1115 165
rect 1117 163 1120 165
rect 1113 161 1120 163
rect 1181 167 1186 170
rect 1188 167 1193 179
rect 1195 167 1203 179
rect 1197 165 1203 167
rect 1197 163 1199 165
rect 1201 163 1203 165
rect 1197 161 1203 163
rect 111 144 118 146
rect 111 142 113 144
rect 115 142 118 144
rect 111 136 118 142
rect 195 144 201 146
rect 195 142 197 144
rect 199 142 201 144
rect 195 140 201 142
rect 226 140 232 142
rect 179 137 184 140
rect 111 134 120 136
rect 100 132 107 134
rect 100 130 102 132
rect 104 130 107 132
rect 100 128 107 130
rect 102 125 107 128
rect 109 125 120 134
rect 122 125 127 136
rect 129 134 136 136
rect 129 132 132 134
rect 134 132 136 134
rect 155 135 164 137
rect 155 133 157 135
rect 159 133 164 135
rect 155 132 164 133
rect 129 130 136 132
rect 129 125 134 130
rect 143 129 148 132
rect 141 127 148 129
rect 141 125 143 127
rect 145 125 148 127
rect 141 123 148 125
rect 150 128 164 132
rect 166 132 174 137
rect 166 130 169 132
rect 171 130 174 132
rect 166 128 174 130
rect 176 134 184 137
rect 176 132 179 134
rect 181 132 184 134
rect 176 128 184 132
rect 186 128 191 140
rect 193 128 201 140
rect 226 138 228 140
rect 230 138 232 140
rect 226 136 232 138
rect 245 140 251 142
rect 266 144 273 146
rect 266 142 268 144
rect 270 142 273 144
rect 245 138 247 140
rect 249 138 251 140
rect 245 136 251 138
rect 226 132 230 136
rect 217 129 222 132
rect 150 123 155 128
rect 215 127 222 129
rect 215 125 217 127
rect 219 125 222 127
rect 215 123 222 125
rect 224 129 230 132
rect 246 129 251 136
rect 266 136 273 142
rect 350 144 356 146
rect 350 142 352 144
rect 354 142 356 144
rect 350 140 356 142
rect 371 144 378 146
rect 371 142 373 144
rect 375 142 378 144
rect 334 137 339 140
rect 266 134 275 136
rect 224 123 232 129
rect 234 127 242 129
rect 234 125 237 127
rect 239 125 242 127
rect 234 123 242 125
rect 244 123 251 129
rect 255 132 262 134
rect 255 130 257 132
rect 259 130 262 132
rect 255 128 262 130
rect 257 125 262 128
rect 264 125 275 134
rect 277 125 282 136
rect 284 134 291 136
rect 284 132 287 134
rect 289 132 291 134
rect 310 135 319 137
rect 310 133 312 135
rect 314 133 319 135
rect 310 132 319 133
rect 284 130 291 132
rect 284 125 289 130
rect 298 129 303 132
rect 296 127 303 129
rect 296 125 298 127
rect 300 125 303 127
rect 296 123 303 125
rect 305 128 319 132
rect 321 132 329 137
rect 321 130 324 132
rect 326 130 329 132
rect 321 128 329 130
rect 331 134 339 137
rect 331 132 334 134
rect 336 132 339 134
rect 331 128 339 132
rect 341 128 346 140
rect 348 128 356 140
rect 371 136 378 142
rect 455 144 461 146
rect 455 142 457 144
rect 459 142 461 144
rect 455 140 461 142
rect 476 140 482 142
rect 439 137 444 140
rect 371 134 380 136
rect 360 132 367 134
rect 360 130 362 132
rect 364 130 367 132
rect 360 128 367 130
rect 305 123 310 128
rect 362 125 367 128
rect 369 125 380 134
rect 382 125 387 136
rect 389 134 396 136
rect 389 132 392 134
rect 394 132 396 134
rect 415 135 424 137
rect 415 133 417 135
rect 419 133 424 135
rect 415 132 424 133
rect 389 130 396 132
rect 389 125 394 130
rect 403 129 408 132
rect 401 127 408 129
rect 401 125 403 127
rect 405 125 408 127
rect 401 123 408 125
rect 410 128 424 132
rect 426 132 434 137
rect 426 130 429 132
rect 431 130 434 132
rect 426 128 434 130
rect 436 134 444 137
rect 436 132 439 134
rect 441 132 444 134
rect 436 128 444 132
rect 446 128 451 140
rect 453 128 461 140
rect 476 138 478 140
rect 480 138 482 140
rect 476 136 482 138
rect 495 140 501 142
rect 516 144 523 146
rect 516 142 518 144
rect 520 142 523 144
rect 495 138 497 140
rect 499 138 501 140
rect 495 136 501 138
rect 476 132 480 136
rect 467 129 472 132
rect 410 123 415 128
rect 465 127 472 129
rect 465 125 467 127
rect 469 125 472 127
rect 465 123 472 125
rect 474 129 480 132
rect 496 129 501 136
rect 516 136 523 142
rect 600 144 606 146
rect 600 142 602 144
rect 604 142 606 144
rect 600 140 606 142
rect 621 144 628 146
rect 621 142 623 144
rect 625 142 628 144
rect 584 137 589 140
rect 516 134 525 136
rect 474 123 482 129
rect 484 127 492 129
rect 484 125 487 127
rect 489 125 492 127
rect 484 123 492 125
rect 494 123 501 129
rect 505 132 512 134
rect 505 130 507 132
rect 509 130 512 132
rect 505 128 512 130
rect 507 125 512 128
rect 514 125 525 134
rect 527 125 532 136
rect 534 134 541 136
rect 534 132 537 134
rect 539 132 541 134
rect 560 135 569 137
rect 560 133 562 135
rect 564 133 569 135
rect 560 132 569 133
rect 534 130 541 132
rect 534 125 539 130
rect 548 129 553 132
rect 546 127 553 129
rect 546 125 548 127
rect 550 125 553 127
rect 546 123 553 125
rect 555 128 569 132
rect 571 132 579 137
rect 571 130 574 132
rect 576 130 579 132
rect 571 128 579 130
rect 581 134 589 137
rect 581 132 584 134
rect 586 132 589 134
rect 581 128 589 132
rect 591 128 596 140
rect 598 128 606 140
rect 621 136 628 142
rect 705 144 711 146
rect 705 142 707 144
rect 709 142 711 144
rect 705 140 711 142
rect 726 140 732 142
rect 689 137 694 140
rect 621 134 630 136
rect 610 132 617 134
rect 610 130 612 132
rect 614 130 617 132
rect 610 128 617 130
rect 555 123 560 128
rect 612 125 617 128
rect 619 125 630 134
rect 632 125 637 136
rect 639 134 646 136
rect 639 132 642 134
rect 644 132 646 134
rect 665 135 674 137
rect 665 133 667 135
rect 669 133 674 135
rect 665 132 674 133
rect 639 130 646 132
rect 639 125 644 130
rect 653 129 658 132
rect 651 127 658 129
rect 651 125 653 127
rect 655 125 658 127
rect 651 123 658 125
rect 660 128 674 132
rect 676 132 684 137
rect 676 130 679 132
rect 681 130 684 132
rect 676 128 684 130
rect 686 134 694 137
rect 686 132 689 134
rect 691 132 694 134
rect 686 128 694 132
rect 696 128 701 140
rect 703 128 711 140
rect 726 138 728 140
rect 730 138 732 140
rect 726 136 732 138
rect 745 140 751 142
rect 766 144 773 146
rect 766 142 768 144
rect 770 142 773 144
rect 745 138 747 140
rect 749 138 751 140
rect 745 136 751 138
rect 726 132 730 136
rect 717 129 722 132
rect 660 123 665 128
rect 715 127 722 129
rect 715 125 717 127
rect 719 125 722 127
rect 715 123 722 125
rect 724 129 730 132
rect 746 129 751 136
rect 766 136 773 142
rect 850 144 856 146
rect 850 142 852 144
rect 854 142 856 144
rect 850 140 856 142
rect 871 144 878 146
rect 871 142 873 144
rect 875 142 878 144
rect 834 137 839 140
rect 766 134 775 136
rect 724 123 732 129
rect 734 127 742 129
rect 734 125 737 127
rect 739 125 742 127
rect 734 123 742 125
rect 744 123 751 129
rect 755 132 762 134
rect 755 130 757 132
rect 759 130 762 132
rect 755 128 762 130
rect 757 125 762 128
rect 764 125 775 134
rect 777 125 782 136
rect 784 134 791 136
rect 784 132 787 134
rect 789 132 791 134
rect 810 135 819 137
rect 810 133 812 135
rect 814 133 819 135
rect 810 132 819 133
rect 784 130 791 132
rect 784 125 789 130
rect 798 129 803 132
rect 796 127 803 129
rect 796 125 798 127
rect 800 125 803 127
rect 796 123 803 125
rect 805 128 819 132
rect 821 132 829 137
rect 821 130 824 132
rect 826 130 829 132
rect 821 128 829 130
rect 831 134 839 137
rect 831 132 834 134
rect 836 132 839 134
rect 831 128 839 132
rect 841 128 846 140
rect 848 128 856 140
rect 871 136 878 142
rect 955 144 961 146
rect 955 142 957 144
rect 959 142 961 144
rect 955 140 961 142
rect 976 140 982 142
rect 939 137 944 140
rect 871 134 880 136
rect 860 132 867 134
rect 860 130 862 132
rect 864 130 867 132
rect 860 128 867 130
rect 805 123 810 128
rect 862 125 867 128
rect 869 125 880 134
rect 882 125 887 136
rect 889 134 896 136
rect 889 132 892 134
rect 894 132 896 134
rect 915 135 924 137
rect 915 133 917 135
rect 919 133 924 135
rect 915 132 924 133
rect 889 130 896 132
rect 889 125 894 130
rect 903 129 908 132
rect 901 127 908 129
rect 901 125 903 127
rect 905 125 908 127
rect 901 123 908 125
rect 910 128 924 132
rect 926 132 934 137
rect 926 130 929 132
rect 931 130 934 132
rect 926 128 934 130
rect 936 134 944 137
rect 936 132 939 134
rect 941 132 944 134
rect 936 128 944 132
rect 946 128 951 140
rect 953 128 961 140
rect 976 138 978 140
rect 980 138 982 140
rect 976 136 982 138
rect 995 140 1001 142
rect 1016 144 1023 146
rect 1016 142 1018 144
rect 1020 142 1023 144
rect 995 138 997 140
rect 999 138 1001 140
rect 995 136 1001 138
rect 976 132 980 136
rect 967 129 972 132
rect 910 123 915 128
rect 965 127 972 129
rect 965 125 967 127
rect 969 125 972 127
rect 965 123 972 125
rect 974 129 980 132
rect 996 129 1001 136
rect 1016 136 1023 142
rect 1100 144 1106 146
rect 1100 142 1102 144
rect 1104 142 1106 144
rect 1100 140 1106 142
rect 1121 144 1128 146
rect 1121 142 1123 144
rect 1125 142 1128 144
rect 1084 137 1089 140
rect 1016 134 1025 136
rect 974 123 982 129
rect 984 127 992 129
rect 984 125 987 127
rect 989 125 992 127
rect 984 123 992 125
rect 994 123 1001 129
rect 1005 132 1012 134
rect 1005 130 1007 132
rect 1009 130 1012 132
rect 1005 128 1012 130
rect 1007 125 1012 128
rect 1014 125 1025 134
rect 1027 125 1032 136
rect 1034 134 1041 136
rect 1034 132 1037 134
rect 1039 132 1041 134
rect 1060 135 1069 137
rect 1060 133 1062 135
rect 1064 133 1069 135
rect 1060 132 1069 133
rect 1034 130 1041 132
rect 1034 125 1039 130
rect 1048 129 1053 132
rect 1046 127 1053 129
rect 1046 125 1048 127
rect 1050 125 1053 127
rect 1046 123 1053 125
rect 1055 128 1069 132
rect 1071 132 1079 137
rect 1071 130 1074 132
rect 1076 130 1079 132
rect 1071 128 1079 130
rect 1081 134 1089 137
rect 1081 132 1084 134
rect 1086 132 1089 134
rect 1081 128 1089 132
rect 1091 128 1096 140
rect 1098 128 1106 140
rect 1121 136 1128 142
rect 1205 144 1211 146
rect 1205 142 1207 144
rect 1209 142 1211 144
rect 1205 140 1211 142
rect 1189 137 1194 140
rect 1121 134 1130 136
rect 1110 132 1117 134
rect 1110 130 1112 132
rect 1114 130 1117 132
rect 1110 128 1117 130
rect 1055 123 1060 128
rect 1112 125 1117 128
rect 1119 125 1130 134
rect 1132 125 1137 136
rect 1139 134 1146 136
rect 1139 132 1142 134
rect 1144 132 1146 134
rect 1165 135 1174 137
rect 1165 133 1167 135
rect 1169 133 1174 135
rect 1165 132 1174 133
rect 1139 130 1146 132
rect 1139 125 1144 130
rect 1153 129 1158 132
rect 1151 127 1158 129
rect 1151 125 1153 127
rect 1155 125 1158 127
rect 1151 123 1158 125
rect 1160 128 1174 132
rect 1176 132 1184 137
rect 1176 130 1179 132
rect 1181 130 1184 132
rect 1176 128 1184 130
rect 1186 134 1194 137
rect 1186 132 1189 134
rect 1191 132 1194 134
rect 1186 128 1194 132
rect 1196 128 1201 140
rect 1203 128 1211 140
rect 1160 123 1165 128
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 9 22 14 25
rect 16 25 24 31
rect 26 29 34 31
rect 26 27 29 29
rect 31 27 34 29
rect 26 25 34 27
rect 36 25 43 31
rect 88 29 95 31
rect 49 26 54 29
rect 16 22 22 25
rect 18 18 22 22
rect 38 18 43 25
rect 47 24 54 26
rect 47 22 49 24
rect 51 22 54 24
rect 47 20 54 22
rect 56 20 67 29
rect 18 16 24 18
rect 18 14 20 16
rect 22 14 24 16
rect 18 12 24 14
rect 37 16 43 18
rect 58 18 67 20
rect 69 18 74 29
rect 76 24 81 29
rect 88 27 90 29
rect 92 27 95 29
rect 88 25 95 27
rect 76 22 83 24
rect 90 22 95 25
rect 97 26 102 31
rect 193 29 200 31
rect 154 26 159 29
rect 97 22 111 26
rect 76 20 79 22
rect 81 20 83 22
rect 76 18 83 20
rect 102 21 111 22
rect 102 19 104 21
rect 106 19 111 21
rect 37 14 39 16
rect 41 14 43 16
rect 37 12 43 14
rect 58 12 65 18
rect 102 17 111 19
rect 113 24 121 26
rect 113 22 116 24
rect 118 22 121 24
rect 113 17 121 22
rect 123 22 131 26
rect 123 20 126 22
rect 128 20 131 22
rect 123 17 131 20
rect 58 10 60 12
rect 62 10 65 12
rect 58 8 65 10
rect 126 14 131 17
rect 133 14 138 26
rect 140 14 148 26
rect 152 24 159 26
rect 152 22 154 24
rect 156 22 159 24
rect 152 20 159 22
rect 161 20 172 29
rect 163 18 172 20
rect 174 18 179 29
rect 181 24 186 29
rect 193 27 195 29
rect 197 27 200 29
rect 193 25 200 27
rect 181 22 188 24
rect 195 22 200 25
rect 202 26 207 31
rect 257 29 264 31
rect 257 27 259 29
rect 261 27 264 29
rect 202 22 216 26
rect 181 20 184 22
rect 186 20 188 22
rect 181 18 188 20
rect 207 21 216 22
rect 207 19 209 21
rect 211 19 216 21
rect 142 12 148 14
rect 142 10 144 12
rect 146 10 148 12
rect 142 8 148 10
rect 163 12 170 18
rect 207 17 216 19
rect 218 24 226 26
rect 218 22 221 24
rect 223 22 226 24
rect 218 17 226 22
rect 228 22 236 26
rect 228 20 231 22
rect 233 20 236 22
rect 228 17 236 20
rect 163 10 165 12
rect 167 10 170 12
rect 163 8 170 10
rect 231 14 236 17
rect 238 14 243 26
rect 245 14 253 26
rect 257 25 264 27
rect 259 22 264 25
rect 266 25 274 31
rect 276 29 284 31
rect 276 27 279 29
rect 281 27 284 29
rect 276 25 284 27
rect 286 25 293 31
rect 338 29 345 31
rect 299 26 304 29
rect 266 22 272 25
rect 268 18 272 22
rect 288 18 293 25
rect 297 24 304 26
rect 297 22 299 24
rect 301 22 304 24
rect 297 20 304 22
rect 306 20 317 29
rect 268 16 274 18
rect 268 14 270 16
rect 272 14 274 16
rect 247 12 253 14
rect 247 10 249 12
rect 251 10 253 12
rect 247 8 253 10
rect 268 12 274 14
rect 287 16 293 18
rect 308 18 317 20
rect 319 18 324 29
rect 326 24 331 29
rect 338 27 340 29
rect 342 27 345 29
rect 338 25 345 27
rect 326 22 333 24
rect 340 22 345 25
rect 347 26 352 31
rect 443 29 450 31
rect 404 26 409 29
rect 347 22 361 26
rect 326 20 329 22
rect 331 20 333 22
rect 326 18 333 20
rect 352 21 361 22
rect 352 19 354 21
rect 356 19 361 21
rect 287 14 289 16
rect 291 14 293 16
rect 287 12 293 14
rect 308 12 315 18
rect 352 17 361 19
rect 363 24 371 26
rect 363 22 366 24
rect 368 22 371 24
rect 363 17 371 22
rect 373 22 381 26
rect 373 20 376 22
rect 378 20 381 22
rect 373 17 381 20
rect 308 10 310 12
rect 312 10 315 12
rect 308 8 315 10
rect 376 14 381 17
rect 383 14 388 26
rect 390 14 398 26
rect 402 24 409 26
rect 402 22 404 24
rect 406 22 409 24
rect 402 20 409 22
rect 411 20 422 29
rect 413 18 422 20
rect 424 18 429 29
rect 431 24 436 29
rect 443 27 445 29
rect 447 27 450 29
rect 443 25 450 27
rect 431 22 438 24
rect 445 22 450 25
rect 452 26 457 31
rect 507 29 514 31
rect 507 27 509 29
rect 511 27 514 29
rect 452 22 466 26
rect 431 20 434 22
rect 436 20 438 22
rect 431 18 438 20
rect 457 21 466 22
rect 457 19 459 21
rect 461 19 466 21
rect 392 12 398 14
rect 392 10 394 12
rect 396 10 398 12
rect 392 8 398 10
rect 413 12 420 18
rect 457 17 466 19
rect 468 24 476 26
rect 468 22 471 24
rect 473 22 476 24
rect 468 17 476 22
rect 478 22 486 26
rect 478 20 481 22
rect 483 20 486 22
rect 478 17 486 20
rect 413 10 415 12
rect 417 10 420 12
rect 413 8 420 10
rect 481 14 486 17
rect 488 14 493 26
rect 495 14 503 26
rect 507 25 514 27
rect 509 22 514 25
rect 516 25 524 31
rect 526 29 534 31
rect 526 27 529 29
rect 531 27 534 29
rect 526 25 534 27
rect 536 25 543 31
rect 588 29 595 31
rect 549 26 554 29
rect 516 22 522 25
rect 518 18 522 22
rect 538 18 543 25
rect 547 24 554 26
rect 547 22 549 24
rect 551 22 554 24
rect 547 20 554 22
rect 556 20 567 29
rect 518 16 524 18
rect 518 14 520 16
rect 522 14 524 16
rect 497 12 503 14
rect 497 10 499 12
rect 501 10 503 12
rect 497 8 503 10
rect 518 12 524 14
rect 537 16 543 18
rect 558 18 567 20
rect 569 18 574 29
rect 576 24 581 29
rect 588 27 590 29
rect 592 27 595 29
rect 588 25 595 27
rect 576 22 583 24
rect 590 22 595 25
rect 597 26 602 31
rect 693 29 700 31
rect 654 26 659 29
rect 597 22 611 26
rect 576 20 579 22
rect 581 20 583 22
rect 576 18 583 20
rect 602 21 611 22
rect 602 19 604 21
rect 606 19 611 21
rect 537 14 539 16
rect 541 14 543 16
rect 537 12 543 14
rect 558 12 565 18
rect 602 17 611 19
rect 613 24 621 26
rect 613 22 616 24
rect 618 22 621 24
rect 613 17 621 22
rect 623 22 631 26
rect 623 20 626 22
rect 628 20 631 22
rect 623 17 631 20
rect 558 10 560 12
rect 562 10 565 12
rect 558 8 565 10
rect 626 14 631 17
rect 633 14 638 26
rect 640 14 648 26
rect 652 24 659 26
rect 652 22 654 24
rect 656 22 659 24
rect 652 20 659 22
rect 661 20 672 29
rect 663 18 672 20
rect 674 18 679 29
rect 681 24 686 29
rect 693 27 695 29
rect 697 27 700 29
rect 693 25 700 27
rect 681 22 688 24
rect 695 22 700 25
rect 702 26 707 31
rect 757 29 764 31
rect 757 27 759 29
rect 761 27 764 29
rect 702 22 716 26
rect 681 20 684 22
rect 686 20 688 22
rect 681 18 688 20
rect 707 21 716 22
rect 707 19 709 21
rect 711 19 716 21
rect 642 12 648 14
rect 642 10 644 12
rect 646 10 648 12
rect 642 8 648 10
rect 663 12 670 18
rect 707 17 716 19
rect 718 24 726 26
rect 718 22 721 24
rect 723 22 726 24
rect 718 17 726 22
rect 728 22 736 26
rect 728 20 731 22
rect 733 20 736 22
rect 728 17 736 20
rect 663 10 665 12
rect 667 10 670 12
rect 663 8 670 10
rect 731 14 736 17
rect 738 14 743 26
rect 745 14 753 26
rect 757 25 764 27
rect 759 22 764 25
rect 766 25 774 31
rect 776 29 784 31
rect 776 27 779 29
rect 781 27 784 29
rect 776 25 784 27
rect 786 25 793 31
rect 838 29 845 31
rect 799 26 804 29
rect 766 22 772 25
rect 768 18 772 22
rect 788 18 793 25
rect 797 24 804 26
rect 797 22 799 24
rect 801 22 804 24
rect 797 20 804 22
rect 806 20 817 29
rect 768 16 774 18
rect 768 14 770 16
rect 772 14 774 16
rect 747 12 753 14
rect 747 10 749 12
rect 751 10 753 12
rect 747 8 753 10
rect 768 12 774 14
rect 787 16 793 18
rect 808 18 817 20
rect 819 18 824 29
rect 826 24 831 29
rect 838 27 840 29
rect 842 27 845 29
rect 838 25 845 27
rect 826 22 833 24
rect 840 22 845 25
rect 847 26 852 31
rect 943 29 950 31
rect 904 26 909 29
rect 847 22 861 26
rect 826 20 829 22
rect 831 20 833 22
rect 826 18 833 20
rect 852 21 861 22
rect 852 19 854 21
rect 856 19 861 21
rect 787 14 789 16
rect 791 14 793 16
rect 787 12 793 14
rect 808 12 815 18
rect 852 17 861 19
rect 863 24 871 26
rect 863 22 866 24
rect 868 22 871 24
rect 863 17 871 22
rect 873 22 881 26
rect 873 20 876 22
rect 878 20 881 22
rect 873 17 881 20
rect 808 10 810 12
rect 812 10 815 12
rect 808 8 815 10
rect 876 14 881 17
rect 883 14 888 26
rect 890 14 898 26
rect 902 24 909 26
rect 902 22 904 24
rect 906 22 909 24
rect 902 20 909 22
rect 911 20 922 29
rect 913 18 922 20
rect 924 18 929 29
rect 931 24 936 29
rect 943 27 945 29
rect 947 27 950 29
rect 943 25 950 27
rect 931 22 938 24
rect 945 22 950 25
rect 952 26 957 31
rect 952 22 966 26
rect 931 20 934 22
rect 936 20 938 22
rect 931 18 938 20
rect 957 21 966 22
rect 957 19 959 21
rect 961 19 966 21
rect 892 12 898 14
rect 892 10 894 12
rect 896 10 898 12
rect 892 8 898 10
rect 913 12 920 18
rect 957 17 966 19
rect 968 24 976 26
rect 968 22 971 24
rect 973 22 976 24
rect 968 17 976 22
rect 978 22 986 26
rect 978 20 981 22
rect 983 20 986 22
rect 978 17 986 20
rect 913 10 915 12
rect 917 10 920 12
rect 913 8 920 10
rect 981 14 986 17
rect 988 14 993 26
rect 995 14 1003 26
rect 997 12 1003 14
rect 997 10 999 12
rect 1001 10 1003 12
rect 997 8 1003 10
<< pdif >>
rect 35 372 41 379
rect 14 363 21 372
rect 14 361 16 363
rect 18 361 21 363
rect 14 359 21 361
rect 23 370 31 372
rect 23 368 26 370
rect 28 368 31 370
rect 23 363 31 368
rect 23 361 26 363
rect 28 361 31 363
rect 23 359 31 361
rect 33 365 41 372
rect 33 363 36 365
rect 38 363 41 365
rect 33 361 41 363
rect 43 377 50 379
rect 43 375 46 377
rect 48 375 50 377
rect 43 370 50 375
rect 75 372 81 379
rect 43 368 46 370
rect 48 368 50 370
rect 43 366 50 368
rect 43 361 48 366
rect 54 363 61 372
rect 54 361 56 363
rect 58 361 61 363
rect 33 359 39 361
rect 54 359 61 361
rect 63 370 71 372
rect 63 368 66 370
rect 68 368 71 370
rect 63 363 71 368
rect 63 361 66 363
rect 68 361 71 363
rect 63 359 71 361
rect 73 365 81 372
rect 73 363 76 365
rect 78 363 81 365
rect 73 361 81 363
rect 83 377 90 379
rect 83 375 86 377
rect 88 375 90 377
rect 83 370 90 375
rect 83 368 86 370
rect 88 368 90 370
rect 83 366 90 368
rect 83 361 88 366
rect 103 364 108 379
rect 101 362 108 364
rect 73 359 79 361
rect 101 360 103 362
rect 105 360 108 362
rect 101 358 108 360
rect 103 352 108 358
rect 110 370 118 379
rect 110 368 113 370
rect 115 368 118 370
rect 110 361 118 368
rect 120 377 128 379
rect 120 375 123 377
rect 125 375 128 377
rect 120 370 128 375
rect 120 368 123 370
rect 125 368 128 370
rect 120 361 128 368
rect 130 363 144 379
rect 130 361 139 363
rect 141 361 144 363
rect 110 352 115 361
rect 132 356 144 361
rect 132 354 139 356
rect 141 354 144 356
rect 132 352 144 354
rect 146 377 153 379
rect 146 375 149 377
rect 151 375 153 377
rect 146 373 153 375
rect 146 352 151 373
rect 187 372 193 379
rect 166 363 173 372
rect 166 361 168 363
rect 170 361 173 363
rect 166 359 173 361
rect 175 370 183 372
rect 175 368 178 370
rect 180 368 183 370
rect 175 363 183 368
rect 175 361 178 363
rect 180 361 183 363
rect 175 359 183 361
rect 185 365 193 372
rect 185 363 188 365
rect 190 363 193 365
rect 185 361 193 363
rect 195 377 202 379
rect 195 375 198 377
rect 200 375 202 377
rect 195 370 202 375
rect 517 374 523 381
rect 195 368 198 370
rect 200 368 202 370
rect 195 366 202 368
rect 195 361 200 366
rect 496 365 503 374
rect 496 363 498 365
rect 500 363 503 365
rect 496 361 503 363
rect 505 372 513 374
rect 505 370 508 372
rect 510 370 513 372
rect 505 365 513 370
rect 505 363 508 365
rect 510 363 513 365
rect 505 361 513 363
rect 515 367 523 374
rect 515 365 518 367
rect 520 365 523 367
rect 515 363 523 365
rect 525 379 532 381
rect 525 377 528 379
rect 530 377 532 379
rect 525 372 532 377
rect 557 374 563 381
rect 525 370 528 372
rect 530 370 532 372
rect 525 368 532 370
rect 525 363 530 368
rect 536 365 543 374
rect 536 363 538 365
rect 540 363 543 365
rect 515 361 521 363
rect 185 359 191 361
rect 536 361 543 363
rect 545 372 553 374
rect 545 370 548 372
rect 550 370 553 372
rect 545 365 553 370
rect 545 363 548 365
rect 550 363 553 365
rect 545 361 553 363
rect 555 367 563 374
rect 555 365 558 367
rect 560 365 563 367
rect 555 363 563 365
rect 565 379 572 381
rect 565 377 568 379
rect 570 377 572 379
rect 565 372 572 377
rect 565 370 568 372
rect 570 370 572 372
rect 565 368 572 370
rect 565 363 570 368
rect 585 366 590 381
rect 583 364 590 366
rect 555 361 561 363
rect 583 362 585 364
rect 587 362 590 364
rect 583 360 590 362
rect 585 354 590 360
rect 592 372 600 381
rect 592 370 595 372
rect 597 370 600 372
rect 592 363 600 370
rect 602 379 610 381
rect 602 377 605 379
rect 607 377 610 379
rect 602 372 610 377
rect 602 370 605 372
rect 607 370 610 372
rect 602 363 610 370
rect 612 365 626 381
rect 612 363 621 365
rect 623 363 626 365
rect 592 354 597 363
rect 614 358 626 363
rect 614 356 621 358
rect 623 356 626 358
rect 614 354 626 356
rect 628 379 635 381
rect 628 377 631 379
rect 633 377 635 379
rect 628 375 635 377
rect 628 354 633 375
rect 669 374 675 381
rect 648 365 655 374
rect 648 363 650 365
rect 652 363 655 365
rect 648 361 655 363
rect 657 372 665 374
rect 657 370 660 372
rect 662 370 665 372
rect 657 365 665 370
rect 657 363 660 365
rect 662 363 665 365
rect 657 361 665 363
rect 667 367 675 374
rect 667 365 670 367
rect 672 365 675 367
rect 667 363 675 365
rect 677 379 684 381
rect 677 377 680 379
rect 682 377 684 379
rect 677 372 684 377
rect 722 374 728 381
rect 677 370 680 372
rect 682 370 684 372
rect 677 368 684 370
rect 677 363 682 368
rect 701 365 708 374
rect 701 363 703 365
rect 705 363 708 365
rect 667 361 673 363
rect 701 361 708 363
rect 710 372 718 374
rect 710 370 713 372
rect 715 370 718 372
rect 710 365 718 370
rect 710 363 713 365
rect 715 363 718 365
rect 710 361 718 363
rect 720 367 728 374
rect 720 365 723 367
rect 725 365 728 367
rect 720 363 728 365
rect 730 379 737 381
rect 730 377 733 379
rect 735 377 737 379
rect 730 372 737 377
rect 762 374 768 381
rect 730 370 733 372
rect 735 370 737 372
rect 730 368 737 370
rect 730 363 735 368
rect 741 365 748 374
rect 741 363 743 365
rect 745 363 748 365
rect 720 361 726 363
rect 741 361 748 363
rect 750 372 758 374
rect 750 370 753 372
rect 755 370 758 372
rect 750 365 758 370
rect 750 363 753 365
rect 755 363 758 365
rect 750 361 758 363
rect 760 367 768 374
rect 760 365 763 367
rect 765 365 768 367
rect 760 363 768 365
rect 770 379 777 381
rect 770 377 773 379
rect 775 377 777 379
rect 770 372 777 377
rect 770 370 773 372
rect 775 370 777 372
rect 770 368 777 370
rect 770 363 775 368
rect 790 366 795 381
rect 788 364 795 366
rect 760 361 766 363
rect 788 362 790 364
rect 792 362 795 364
rect 788 360 795 362
rect 790 354 795 360
rect 797 372 805 381
rect 797 370 800 372
rect 802 370 805 372
rect 797 363 805 370
rect 807 379 815 381
rect 807 377 810 379
rect 812 377 815 379
rect 807 372 815 377
rect 807 370 810 372
rect 812 370 815 372
rect 807 363 815 370
rect 817 365 831 381
rect 817 363 826 365
rect 828 363 831 365
rect 797 354 802 363
rect 819 358 831 363
rect 819 356 826 358
rect 828 356 831 358
rect 819 354 831 356
rect 833 379 840 381
rect 833 377 836 379
rect 838 377 840 379
rect 833 375 840 377
rect 833 354 838 375
rect 874 374 880 381
rect 853 365 860 374
rect 853 363 855 365
rect 857 363 860 365
rect 853 361 860 363
rect 862 372 870 374
rect 862 370 865 372
rect 867 370 870 372
rect 862 365 870 370
rect 862 363 865 365
rect 867 363 870 365
rect 862 361 870 363
rect 872 367 880 374
rect 872 365 875 367
rect 877 365 880 367
rect 872 363 880 365
rect 882 379 889 381
rect 882 377 885 379
rect 887 377 889 379
rect 882 372 889 377
rect 882 370 885 372
rect 887 370 889 372
rect 882 368 889 370
rect 882 363 887 368
rect 872 361 878 363
rect 25 331 31 333
rect 16 326 21 331
rect 14 324 21 326
rect 14 322 16 324
rect 18 322 21 324
rect 14 317 21 322
rect 14 315 16 317
rect 18 315 21 317
rect 14 313 21 315
rect 23 329 31 331
rect 23 327 26 329
rect 28 327 31 329
rect 23 320 31 327
rect 33 331 41 333
rect 33 329 36 331
rect 38 329 41 331
rect 33 324 41 329
rect 33 322 36 324
rect 38 322 41 324
rect 33 320 41 322
rect 43 331 50 333
rect 43 329 46 331
rect 48 329 50 331
rect 43 320 50 329
rect 54 331 61 333
rect 54 329 56 331
rect 58 329 61 331
rect 54 320 61 329
rect 63 331 71 333
rect 63 329 66 331
rect 68 329 71 331
rect 63 324 71 329
rect 63 322 66 324
rect 68 322 71 324
rect 63 320 71 322
rect 73 331 79 333
rect 105 331 111 333
rect 73 329 81 331
rect 73 327 76 329
rect 78 327 81 329
rect 73 320 81 327
rect 23 313 29 320
rect 75 313 81 320
rect 83 326 88 331
rect 96 326 101 331
rect 83 324 90 326
rect 83 322 86 324
rect 88 322 90 324
rect 83 317 90 322
rect 83 315 86 317
rect 88 315 90 317
rect 83 313 90 315
rect 94 324 101 326
rect 94 322 96 324
rect 98 322 101 324
rect 94 317 101 322
rect 94 315 96 317
rect 98 315 101 317
rect 94 313 101 315
rect 103 329 111 331
rect 103 327 106 329
rect 108 327 111 329
rect 103 320 111 327
rect 113 331 121 333
rect 113 329 116 331
rect 118 329 121 331
rect 113 324 121 329
rect 113 322 116 324
rect 118 322 121 324
rect 113 320 121 322
rect 123 331 130 333
rect 123 329 126 331
rect 128 329 130 331
rect 123 320 130 329
rect 103 313 109 320
rect 145 319 150 340
rect 143 317 150 319
rect 143 315 145 317
rect 147 315 150 317
rect 143 313 150 315
rect 152 338 164 340
rect 152 336 155 338
rect 157 336 164 338
rect 152 331 164 336
rect 181 331 186 340
rect 152 329 155 331
rect 157 329 166 331
rect 152 313 166 329
rect 168 324 176 331
rect 168 322 171 324
rect 173 322 176 324
rect 168 317 176 322
rect 168 315 171 317
rect 173 315 176 317
rect 168 313 176 315
rect 178 324 186 331
rect 178 322 181 324
rect 183 322 186 324
rect 178 313 186 322
rect 188 334 193 340
rect 188 332 195 334
rect 507 333 513 335
rect 188 330 191 332
rect 193 330 195 332
rect 188 328 195 330
rect 498 328 503 333
rect 188 313 193 328
rect 496 326 503 328
rect 496 324 498 326
rect 500 324 503 326
rect 496 319 503 324
rect 496 317 498 319
rect 500 317 503 319
rect 496 315 503 317
rect 505 331 513 333
rect 505 329 508 331
rect 510 329 513 331
rect 505 322 513 329
rect 515 333 523 335
rect 515 331 518 333
rect 520 331 523 333
rect 515 326 523 331
rect 515 324 518 326
rect 520 324 523 326
rect 515 322 523 324
rect 525 333 532 335
rect 525 331 528 333
rect 530 331 532 333
rect 525 322 532 331
rect 536 333 543 335
rect 536 331 538 333
rect 540 331 543 333
rect 536 322 543 331
rect 545 333 553 335
rect 545 331 548 333
rect 550 331 553 333
rect 545 326 553 331
rect 545 324 548 326
rect 550 324 553 326
rect 545 322 553 324
rect 555 333 561 335
rect 587 333 593 335
rect 555 331 563 333
rect 555 329 558 331
rect 560 329 563 331
rect 555 322 563 329
rect 505 315 511 322
rect 557 315 563 322
rect 565 328 570 333
rect 578 328 583 333
rect 565 326 572 328
rect 565 324 568 326
rect 570 324 572 326
rect 565 319 572 324
rect 565 317 568 319
rect 570 317 572 319
rect 565 315 572 317
rect 576 326 583 328
rect 576 324 578 326
rect 580 324 583 326
rect 576 319 583 324
rect 576 317 578 319
rect 580 317 583 319
rect 576 315 583 317
rect 585 331 593 333
rect 585 329 588 331
rect 590 329 593 331
rect 585 322 593 329
rect 595 333 603 335
rect 595 331 598 333
rect 600 331 603 333
rect 595 326 603 331
rect 595 324 598 326
rect 600 324 603 326
rect 595 322 603 324
rect 605 333 612 335
rect 605 331 608 333
rect 610 331 612 333
rect 605 322 612 331
rect 585 315 591 322
rect 627 321 632 342
rect 625 319 632 321
rect 625 317 627 319
rect 629 317 632 319
rect 625 315 632 317
rect 634 340 646 342
rect 634 338 637 340
rect 639 338 646 340
rect 634 333 646 338
rect 663 333 668 342
rect 634 331 637 333
rect 639 331 648 333
rect 634 315 648 331
rect 650 326 658 333
rect 650 324 653 326
rect 655 324 658 326
rect 650 319 658 324
rect 650 317 653 319
rect 655 317 658 319
rect 650 315 658 317
rect 660 326 668 333
rect 660 324 663 326
rect 665 324 668 326
rect 660 315 668 324
rect 670 336 675 342
rect 670 334 677 336
rect 670 332 673 334
rect 675 332 677 334
rect 712 333 718 335
rect 670 330 677 332
rect 670 315 675 330
rect 703 328 708 333
rect 701 326 708 328
rect 701 324 703 326
rect 705 324 708 326
rect 701 319 708 324
rect 701 317 703 319
rect 705 317 708 319
rect 701 315 708 317
rect 710 331 718 333
rect 710 329 713 331
rect 715 329 718 331
rect 710 322 718 329
rect 720 333 728 335
rect 720 331 723 333
rect 725 331 728 333
rect 720 326 728 331
rect 720 324 723 326
rect 725 324 728 326
rect 720 322 728 324
rect 730 333 737 335
rect 730 331 733 333
rect 735 331 737 333
rect 730 322 737 331
rect 741 333 748 335
rect 741 331 743 333
rect 745 331 748 333
rect 741 322 748 331
rect 750 333 758 335
rect 750 331 753 333
rect 755 331 758 333
rect 750 326 758 331
rect 750 324 753 326
rect 755 324 758 326
rect 750 322 758 324
rect 760 333 766 335
rect 792 333 798 335
rect 760 331 768 333
rect 760 329 763 331
rect 765 329 768 331
rect 760 322 768 329
rect 710 315 716 322
rect 762 315 768 322
rect 770 328 775 333
rect 783 328 788 333
rect 770 326 777 328
rect 770 324 773 326
rect 775 324 777 326
rect 770 319 777 324
rect 770 317 773 319
rect 775 317 777 319
rect 770 315 777 317
rect 781 326 788 328
rect 781 324 783 326
rect 785 324 788 326
rect 781 319 788 324
rect 781 317 783 319
rect 785 317 788 319
rect 781 315 788 317
rect 790 331 798 333
rect 790 329 793 331
rect 795 329 798 331
rect 790 322 798 329
rect 800 333 808 335
rect 800 331 803 333
rect 805 331 808 333
rect 800 326 808 331
rect 800 324 803 326
rect 805 324 808 326
rect 800 322 808 324
rect 810 333 817 335
rect 810 331 813 333
rect 815 331 817 333
rect 810 322 817 331
rect 790 315 796 322
rect 832 321 837 342
rect 830 319 837 321
rect 830 317 832 319
rect 834 317 837 319
rect 830 315 837 317
rect 839 340 851 342
rect 839 338 842 340
rect 844 338 851 340
rect 839 333 851 338
rect 868 333 873 342
rect 839 331 842 333
rect 844 331 853 333
rect 839 315 853 331
rect 855 326 863 333
rect 855 324 858 326
rect 860 324 863 326
rect 855 319 863 324
rect 855 317 858 319
rect 860 317 863 319
rect 855 315 863 317
rect 865 326 873 333
rect 865 324 868 326
rect 870 324 873 326
rect 865 315 873 324
rect 875 336 880 342
rect 875 334 882 336
rect 875 332 878 334
rect 880 332 882 334
rect 875 330 882 332
rect 875 315 880 330
rect 1043 256 1049 263
rect 1022 247 1029 256
rect 1022 245 1024 247
rect 1026 245 1029 247
rect 1022 243 1029 245
rect 1031 254 1039 256
rect 1031 252 1034 254
rect 1036 252 1039 254
rect 1031 247 1039 252
rect 1031 245 1034 247
rect 1036 245 1039 247
rect 1031 243 1039 245
rect 1041 249 1049 256
rect 1041 247 1044 249
rect 1046 247 1049 249
rect 1041 245 1049 247
rect 1051 261 1058 263
rect 1051 259 1054 261
rect 1056 259 1058 261
rect 1051 254 1058 259
rect 1083 256 1089 263
rect 1051 252 1054 254
rect 1056 252 1058 254
rect 1051 250 1058 252
rect 1051 245 1056 250
rect 1062 247 1069 256
rect 1062 245 1064 247
rect 1066 245 1069 247
rect 1041 243 1047 245
rect 1062 243 1069 245
rect 1071 254 1079 256
rect 1071 252 1074 254
rect 1076 252 1079 254
rect 1071 247 1079 252
rect 1071 245 1074 247
rect 1076 245 1079 247
rect 1071 243 1079 245
rect 1081 249 1089 256
rect 1081 247 1084 249
rect 1086 247 1089 249
rect 1081 245 1089 247
rect 1091 261 1098 263
rect 1091 259 1094 261
rect 1096 259 1098 261
rect 1091 254 1098 259
rect 1091 252 1094 254
rect 1096 252 1098 254
rect 1091 250 1098 252
rect 1091 245 1096 250
rect 1111 248 1116 263
rect 1109 246 1116 248
rect 1081 243 1087 245
rect 1109 244 1111 246
rect 1113 244 1116 246
rect 1109 242 1116 244
rect 1111 236 1116 242
rect 1118 254 1126 263
rect 1118 252 1121 254
rect 1123 252 1126 254
rect 1118 245 1126 252
rect 1128 261 1136 263
rect 1128 259 1131 261
rect 1133 259 1136 261
rect 1128 254 1136 259
rect 1128 252 1131 254
rect 1133 252 1136 254
rect 1128 245 1136 252
rect 1138 247 1152 263
rect 1138 245 1147 247
rect 1149 245 1152 247
rect 1118 236 1123 245
rect 1140 240 1152 245
rect 1140 238 1147 240
rect 1149 238 1152 240
rect 1140 236 1152 238
rect 1154 261 1161 263
rect 1154 259 1157 261
rect 1159 259 1161 261
rect 1154 257 1161 259
rect 1154 236 1159 257
rect 1195 256 1201 263
rect 1174 247 1181 256
rect 1174 245 1176 247
rect 1178 245 1181 247
rect 1174 243 1181 245
rect 1183 254 1191 256
rect 1183 252 1186 254
rect 1188 252 1191 254
rect 1183 247 1191 252
rect 1183 245 1186 247
rect 1188 245 1191 247
rect 1183 243 1191 245
rect 1193 249 1201 256
rect 1193 247 1196 249
rect 1198 247 1201 249
rect 1193 245 1201 247
rect 1203 261 1210 263
rect 1203 259 1206 261
rect 1208 259 1210 261
rect 1203 254 1210 259
rect 1203 252 1206 254
rect 1208 252 1210 254
rect 1203 250 1210 252
rect 1203 245 1208 250
rect 1193 243 1199 245
rect 12 222 21 224
rect 12 220 14 222
rect 16 220 21 222
rect 12 214 21 220
rect 1 212 8 214
rect 1 210 3 212
rect 5 210 8 212
rect 1 205 8 210
rect 1 203 3 205
rect 5 203 8 205
rect 1 201 8 203
rect 3 196 8 201
rect 10 203 21 214
rect 23 203 28 224
rect 30 217 35 224
rect 30 215 37 217
rect 52 215 58 217
rect 30 213 33 215
rect 35 213 37 215
rect 30 211 37 213
rect 30 203 35 211
rect 43 210 48 215
rect 41 208 48 210
rect 41 206 43 208
rect 45 206 48 208
rect 10 196 18 203
rect 41 201 48 206
rect 41 199 43 201
rect 45 199 48 201
rect 41 197 48 199
rect 50 213 58 215
rect 50 211 53 213
rect 55 211 58 213
rect 50 204 58 211
rect 60 215 68 217
rect 60 213 63 215
rect 65 213 68 215
rect 60 208 68 213
rect 60 206 63 208
rect 65 206 68 208
rect 60 204 68 206
rect 70 215 77 217
rect 70 213 73 215
rect 75 213 77 215
rect 70 204 77 213
rect 50 197 56 204
rect 92 203 97 224
rect 90 201 97 203
rect 90 199 92 201
rect 94 199 97 201
rect 90 197 97 199
rect 99 222 111 224
rect 99 220 102 222
rect 104 220 111 222
rect 99 215 111 220
rect 128 215 133 224
rect 99 213 102 215
rect 104 213 113 215
rect 99 197 113 213
rect 115 208 123 215
rect 115 206 118 208
rect 120 206 123 208
rect 115 201 123 206
rect 115 199 118 201
rect 120 199 123 201
rect 115 197 123 199
rect 125 208 133 215
rect 125 206 128 208
rect 130 206 133 208
rect 125 197 133 206
rect 135 218 140 224
rect 135 216 142 218
rect 135 214 138 216
rect 140 214 142 216
rect 157 215 163 217
rect 135 212 142 214
rect 135 197 140 212
rect 148 210 153 215
rect 146 208 153 210
rect 146 206 148 208
rect 150 206 153 208
rect 146 201 153 206
rect 146 199 148 201
rect 150 199 153 201
rect 146 197 153 199
rect 155 213 163 215
rect 155 211 158 213
rect 160 211 163 213
rect 155 204 163 211
rect 165 215 173 217
rect 165 213 168 215
rect 170 213 173 215
rect 165 208 173 213
rect 165 206 168 208
rect 170 206 173 208
rect 165 204 173 206
rect 175 215 182 217
rect 175 213 178 215
rect 180 213 182 215
rect 175 204 182 213
rect 155 197 161 204
rect 197 203 202 224
rect 195 201 202 203
rect 195 199 197 201
rect 199 199 202 201
rect 195 197 202 199
rect 204 222 216 224
rect 204 220 207 222
rect 209 220 216 222
rect 204 215 216 220
rect 233 215 238 224
rect 204 213 207 215
rect 209 213 218 215
rect 204 197 218 213
rect 220 208 228 215
rect 220 206 223 208
rect 225 206 228 208
rect 220 201 228 206
rect 220 199 223 201
rect 225 199 228 201
rect 220 197 228 199
rect 230 208 238 215
rect 230 206 233 208
rect 235 206 238 208
rect 230 197 238 206
rect 240 218 245 224
rect 262 222 271 224
rect 262 220 264 222
rect 266 220 271 222
rect 240 216 247 218
rect 240 214 243 216
rect 245 214 247 216
rect 262 214 271 220
rect 240 212 247 214
rect 251 212 258 214
rect 240 197 245 212
rect 251 210 253 212
rect 255 210 258 212
rect 251 205 258 210
rect 251 203 253 205
rect 255 203 258 205
rect 251 201 258 203
rect 253 196 258 201
rect 260 203 271 214
rect 273 203 278 224
rect 280 217 285 224
rect 280 215 287 217
rect 302 215 308 217
rect 280 213 283 215
rect 285 213 287 215
rect 280 211 287 213
rect 280 203 285 211
rect 293 210 298 215
rect 291 208 298 210
rect 291 206 293 208
rect 295 206 298 208
rect 260 196 268 203
rect 291 201 298 206
rect 291 199 293 201
rect 295 199 298 201
rect 291 197 298 199
rect 300 213 308 215
rect 300 211 303 213
rect 305 211 308 213
rect 300 204 308 211
rect 310 215 318 217
rect 310 213 313 215
rect 315 213 318 215
rect 310 208 318 213
rect 310 206 313 208
rect 315 206 318 208
rect 310 204 318 206
rect 320 215 327 217
rect 320 213 323 215
rect 325 213 327 215
rect 320 204 327 213
rect 300 197 306 204
rect 342 203 347 224
rect 340 201 347 203
rect 340 199 342 201
rect 344 199 347 201
rect 340 197 347 199
rect 349 222 361 224
rect 349 220 352 222
rect 354 220 361 222
rect 349 215 361 220
rect 378 215 383 224
rect 349 213 352 215
rect 354 213 363 215
rect 349 197 363 213
rect 365 208 373 215
rect 365 206 368 208
rect 370 206 373 208
rect 365 201 373 206
rect 365 199 368 201
rect 370 199 373 201
rect 365 197 373 199
rect 375 208 383 215
rect 375 206 378 208
rect 380 206 383 208
rect 375 197 383 206
rect 385 218 390 224
rect 385 216 392 218
rect 385 214 388 216
rect 390 214 392 216
rect 407 215 413 217
rect 385 212 392 214
rect 385 197 390 212
rect 398 210 403 215
rect 396 208 403 210
rect 396 206 398 208
rect 400 206 403 208
rect 396 201 403 206
rect 396 199 398 201
rect 400 199 403 201
rect 396 197 403 199
rect 405 213 413 215
rect 405 211 408 213
rect 410 211 413 213
rect 405 204 413 211
rect 415 215 423 217
rect 415 213 418 215
rect 420 213 423 215
rect 415 208 423 213
rect 415 206 418 208
rect 420 206 423 208
rect 415 204 423 206
rect 425 215 432 217
rect 425 213 428 215
rect 430 213 432 215
rect 425 204 432 213
rect 405 197 411 204
rect 447 203 452 224
rect 445 201 452 203
rect 445 199 447 201
rect 449 199 452 201
rect 445 197 452 199
rect 454 222 466 224
rect 454 220 457 222
rect 459 220 466 222
rect 454 215 466 220
rect 483 215 488 224
rect 454 213 457 215
rect 459 213 468 215
rect 454 197 468 213
rect 470 208 478 215
rect 470 206 473 208
rect 475 206 478 208
rect 470 201 478 206
rect 470 199 473 201
rect 475 199 478 201
rect 470 197 478 199
rect 480 208 488 215
rect 480 206 483 208
rect 485 206 488 208
rect 480 197 488 206
rect 490 218 495 224
rect 512 222 521 224
rect 512 220 514 222
rect 516 220 521 222
rect 490 216 497 218
rect 490 214 493 216
rect 495 214 497 216
rect 512 214 521 220
rect 490 212 497 214
rect 501 212 508 214
rect 490 197 495 212
rect 501 210 503 212
rect 505 210 508 212
rect 501 205 508 210
rect 501 203 503 205
rect 505 203 508 205
rect 501 201 508 203
rect 503 196 508 201
rect 510 203 521 214
rect 523 203 528 224
rect 530 217 535 224
rect 530 215 537 217
rect 552 215 558 217
rect 530 213 533 215
rect 535 213 537 215
rect 530 211 537 213
rect 530 203 535 211
rect 543 210 548 215
rect 541 208 548 210
rect 541 206 543 208
rect 545 206 548 208
rect 510 196 518 203
rect 541 201 548 206
rect 541 199 543 201
rect 545 199 548 201
rect 541 197 548 199
rect 550 213 558 215
rect 550 211 553 213
rect 555 211 558 213
rect 550 204 558 211
rect 560 215 568 217
rect 560 213 563 215
rect 565 213 568 215
rect 560 208 568 213
rect 560 206 563 208
rect 565 206 568 208
rect 560 204 568 206
rect 570 215 577 217
rect 570 213 573 215
rect 575 213 577 215
rect 570 204 577 213
rect 550 197 556 204
rect 592 203 597 224
rect 590 201 597 203
rect 590 199 592 201
rect 594 199 597 201
rect 590 197 597 199
rect 599 222 611 224
rect 599 220 602 222
rect 604 220 611 222
rect 599 215 611 220
rect 628 215 633 224
rect 599 213 602 215
rect 604 213 613 215
rect 599 197 613 213
rect 615 208 623 215
rect 615 206 618 208
rect 620 206 623 208
rect 615 201 623 206
rect 615 199 618 201
rect 620 199 623 201
rect 615 197 623 199
rect 625 208 633 215
rect 625 206 628 208
rect 630 206 633 208
rect 625 197 633 206
rect 635 218 640 224
rect 635 216 642 218
rect 635 214 638 216
rect 640 214 642 216
rect 657 215 663 217
rect 635 212 642 214
rect 635 197 640 212
rect 648 210 653 215
rect 646 208 653 210
rect 646 206 648 208
rect 650 206 653 208
rect 646 201 653 206
rect 646 199 648 201
rect 650 199 653 201
rect 646 197 653 199
rect 655 213 663 215
rect 655 211 658 213
rect 660 211 663 213
rect 655 204 663 211
rect 665 215 673 217
rect 665 213 668 215
rect 670 213 673 215
rect 665 208 673 213
rect 665 206 668 208
rect 670 206 673 208
rect 665 204 673 206
rect 675 215 682 217
rect 675 213 678 215
rect 680 213 682 215
rect 675 204 682 213
rect 655 197 661 204
rect 697 203 702 224
rect 695 201 702 203
rect 695 199 697 201
rect 699 199 702 201
rect 695 197 702 199
rect 704 222 716 224
rect 704 220 707 222
rect 709 220 716 222
rect 704 215 716 220
rect 733 215 738 224
rect 704 213 707 215
rect 709 213 718 215
rect 704 197 718 213
rect 720 208 728 215
rect 720 206 723 208
rect 725 206 728 208
rect 720 201 728 206
rect 720 199 723 201
rect 725 199 728 201
rect 720 197 728 199
rect 730 208 738 215
rect 730 206 733 208
rect 735 206 738 208
rect 730 197 738 206
rect 740 218 745 224
rect 762 222 771 224
rect 762 220 764 222
rect 766 220 771 222
rect 740 216 747 218
rect 740 214 743 216
rect 745 214 747 216
rect 762 214 771 220
rect 740 212 747 214
rect 751 212 758 214
rect 740 197 745 212
rect 751 210 753 212
rect 755 210 758 212
rect 751 205 758 210
rect 751 203 753 205
rect 755 203 758 205
rect 751 201 758 203
rect 753 196 758 201
rect 760 203 771 214
rect 773 203 778 224
rect 780 217 785 224
rect 780 215 787 217
rect 802 215 808 217
rect 780 213 783 215
rect 785 213 787 215
rect 780 211 787 213
rect 780 203 785 211
rect 793 210 798 215
rect 791 208 798 210
rect 791 206 793 208
rect 795 206 798 208
rect 760 196 768 203
rect 791 201 798 206
rect 791 199 793 201
rect 795 199 798 201
rect 791 197 798 199
rect 800 213 808 215
rect 800 211 803 213
rect 805 211 808 213
rect 800 204 808 211
rect 810 215 818 217
rect 810 213 813 215
rect 815 213 818 215
rect 810 208 818 213
rect 810 206 813 208
rect 815 206 818 208
rect 810 204 818 206
rect 820 215 827 217
rect 820 213 823 215
rect 825 213 827 215
rect 820 204 827 213
rect 800 197 806 204
rect 842 203 847 224
rect 840 201 847 203
rect 840 199 842 201
rect 844 199 847 201
rect 840 197 847 199
rect 849 222 861 224
rect 849 220 852 222
rect 854 220 861 222
rect 849 215 861 220
rect 878 215 883 224
rect 849 213 852 215
rect 854 213 863 215
rect 849 197 863 213
rect 865 208 873 215
rect 865 206 868 208
rect 870 206 873 208
rect 865 201 873 206
rect 865 199 868 201
rect 870 199 873 201
rect 865 197 873 199
rect 875 208 883 215
rect 875 206 878 208
rect 880 206 883 208
rect 875 197 883 206
rect 885 218 890 224
rect 885 216 892 218
rect 885 214 888 216
rect 890 214 892 216
rect 907 215 913 217
rect 885 212 892 214
rect 885 197 890 212
rect 898 210 903 215
rect 896 208 903 210
rect 896 206 898 208
rect 900 206 903 208
rect 896 201 903 206
rect 896 199 898 201
rect 900 199 903 201
rect 896 197 903 199
rect 905 213 913 215
rect 905 211 908 213
rect 910 211 913 213
rect 905 204 913 211
rect 915 215 923 217
rect 915 213 918 215
rect 920 213 923 215
rect 915 208 923 213
rect 915 206 918 208
rect 920 206 923 208
rect 915 204 923 206
rect 925 215 932 217
rect 925 213 928 215
rect 930 213 932 215
rect 925 204 932 213
rect 905 197 911 204
rect 947 203 952 224
rect 945 201 952 203
rect 945 199 947 201
rect 949 199 952 201
rect 945 197 952 199
rect 954 222 966 224
rect 954 220 957 222
rect 959 220 966 222
rect 954 215 966 220
rect 983 215 988 224
rect 954 213 957 215
rect 959 213 968 215
rect 954 197 968 213
rect 970 208 978 215
rect 970 206 973 208
rect 975 206 978 208
rect 970 201 978 206
rect 970 199 973 201
rect 975 199 978 201
rect 970 197 978 199
rect 980 208 988 215
rect 980 206 983 208
rect 985 206 988 208
rect 980 197 988 206
rect 990 218 995 224
rect 990 216 997 218
rect 990 214 993 216
rect 995 214 997 216
rect 1033 215 1039 217
rect 990 212 997 214
rect 990 197 995 212
rect 1024 210 1029 215
rect 1022 208 1029 210
rect 1022 206 1024 208
rect 1026 206 1029 208
rect 1022 201 1029 206
rect 1022 199 1024 201
rect 1026 199 1029 201
rect 1022 197 1029 199
rect 1031 213 1039 215
rect 1031 211 1034 213
rect 1036 211 1039 213
rect 1031 204 1039 211
rect 1041 215 1049 217
rect 1041 213 1044 215
rect 1046 213 1049 215
rect 1041 208 1049 213
rect 1041 206 1044 208
rect 1046 206 1049 208
rect 1041 204 1049 206
rect 1051 215 1058 217
rect 1051 213 1054 215
rect 1056 213 1058 215
rect 1051 204 1058 213
rect 1062 215 1069 217
rect 1062 213 1064 215
rect 1066 213 1069 215
rect 1062 204 1069 213
rect 1071 215 1079 217
rect 1071 213 1074 215
rect 1076 213 1079 215
rect 1071 208 1079 213
rect 1071 206 1074 208
rect 1076 206 1079 208
rect 1071 204 1079 206
rect 1081 215 1087 217
rect 1113 215 1119 217
rect 1081 213 1089 215
rect 1081 211 1084 213
rect 1086 211 1089 213
rect 1081 204 1089 211
rect 1031 197 1037 204
rect 1083 197 1089 204
rect 1091 210 1096 215
rect 1104 210 1109 215
rect 1091 208 1098 210
rect 1091 206 1094 208
rect 1096 206 1098 208
rect 1091 201 1098 206
rect 1091 199 1094 201
rect 1096 199 1098 201
rect 1091 197 1098 199
rect 1102 208 1109 210
rect 1102 206 1104 208
rect 1106 206 1109 208
rect 1102 201 1109 206
rect 1102 199 1104 201
rect 1106 199 1109 201
rect 1102 197 1109 199
rect 1111 213 1119 215
rect 1111 211 1114 213
rect 1116 211 1119 213
rect 1111 204 1119 211
rect 1121 215 1129 217
rect 1121 213 1124 215
rect 1126 213 1129 215
rect 1121 208 1129 213
rect 1121 206 1124 208
rect 1126 206 1129 208
rect 1121 204 1129 206
rect 1131 215 1138 217
rect 1131 213 1134 215
rect 1136 213 1138 215
rect 1131 204 1138 213
rect 1111 197 1117 204
rect 1153 203 1158 224
rect 1151 201 1158 203
rect 1151 199 1153 201
rect 1155 199 1158 201
rect 1151 197 1158 199
rect 1160 222 1172 224
rect 1160 220 1163 222
rect 1165 220 1172 222
rect 1160 215 1172 220
rect 1189 215 1194 224
rect 1160 213 1163 215
rect 1165 213 1174 215
rect 1160 197 1174 213
rect 1176 208 1184 215
rect 1176 206 1179 208
rect 1181 206 1184 208
rect 1176 201 1184 206
rect 1176 199 1179 201
rect 1181 199 1184 201
rect 1176 197 1184 199
rect 1186 208 1194 215
rect 1186 206 1189 208
rect 1191 206 1194 208
rect 1186 197 1194 206
rect 1196 218 1201 224
rect 1196 216 1203 218
rect 1196 214 1199 216
rect 1201 214 1203 216
rect 1196 212 1203 214
rect 1196 197 1201 212
rect 100 108 107 110
rect 100 106 102 108
rect 104 106 107 108
rect 100 101 107 106
rect 100 99 102 101
rect 104 99 107 101
rect 100 97 107 99
rect 102 92 107 97
rect 109 103 115 110
rect 149 108 156 110
rect 149 106 151 108
rect 153 106 156 108
rect 149 104 156 106
rect 109 96 117 103
rect 109 94 112 96
rect 114 94 117 96
rect 109 92 117 94
rect 111 90 117 92
rect 119 101 127 103
rect 119 99 122 101
rect 124 99 127 101
rect 119 94 127 99
rect 119 92 122 94
rect 124 92 127 94
rect 119 90 127 92
rect 129 94 136 103
rect 129 92 132 94
rect 134 92 136 94
rect 129 90 136 92
rect 151 83 156 104
rect 158 94 172 110
rect 158 92 161 94
rect 163 92 172 94
rect 174 108 182 110
rect 174 106 177 108
rect 179 106 182 108
rect 174 101 182 106
rect 174 99 177 101
rect 179 99 182 101
rect 174 92 182 99
rect 184 101 192 110
rect 184 99 187 101
rect 189 99 192 101
rect 184 92 192 99
rect 158 87 170 92
rect 158 85 161 87
rect 163 85 170 87
rect 158 83 170 85
rect 187 83 192 92
rect 194 95 199 110
rect 217 106 222 111
rect 215 104 222 106
rect 215 102 217 104
rect 219 102 222 104
rect 215 97 222 102
rect 215 95 217 97
rect 219 95 222 97
rect 194 93 201 95
rect 215 93 222 95
rect 224 104 232 111
rect 255 108 262 110
rect 255 106 257 108
rect 259 106 262 108
rect 224 93 235 104
rect 194 91 197 93
rect 199 91 201 93
rect 194 89 201 91
rect 194 83 199 89
rect 226 87 235 93
rect 226 85 228 87
rect 230 85 235 87
rect 226 83 235 85
rect 237 83 242 104
rect 244 96 249 104
rect 255 101 262 106
rect 255 99 257 101
rect 259 99 262 101
rect 255 97 262 99
rect 244 94 251 96
rect 244 92 247 94
rect 249 92 251 94
rect 257 92 262 97
rect 264 103 270 110
rect 304 108 311 110
rect 304 106 306 108
rect 308 106 311 108
rect 304 104 311 106
rect 264 96 272 103
rect 264 94 267 96
rect 269 94 272 96
rect 264 92 272 94
rect 244 90 251 92
rect 244 83 249 90
rect 266 90 272 92
rect 274 101 282 103
rect 274 99 277 101
rect 279 99 282 101
rect 274 94 282 99
rect 274 92 277 94
rect 279 92 282 94
rect 274 90 282 92
rect 284 94 291 103
rect 284 92 287 94
rect 289 92 291 94
rect 284 90 291 92
rect 306 83 311 104
rect 313 94 327 110
rect 313 92 316 94
rect 318 92 327 94
rect 329 108 337 110
rect 329 106 332 108
rect 334 106 337 108
rect 329 101 337 106
rect 329 99 332 101
rect 334 99 337 101
rect 329 92 337 99
rect 339 101 347 110
rect 339 99 342 101
rect 344 99 347 101
rect 339 92 347 99
rect 313 87 325 92
rect 313 85 316 87
rect 318 85 325 87
rect 313 83 325 85
rect 342 83 347 92
rect 349 95 354 110
rect 360 108 367 110
rect 360 106 362 108
rect 364 106 367 108
rect 360 101 367 106
rect 360 99 362 101
rect 364 99 367 101
rect 360 97 367 99
rect 349 93 356 95
rect 349 91 352 93
rect 354 91 356 93
rect 362 92 367 97
rect 369 103 375 110
rect 409 108 416 110
rect 409 106 411 108
rect 413 106 416 108
rect 409 104 416 106
rect 369 96 377 103
rect 369 94 372 96
rect 374 94 377 96
rect 369 92 377 94
rect 349 89 356 91
rect 349 83 354 89
rect 371 90 377 92
rect 379 101 387 103
rect 379 99 382 101
rect 384 99 387 101
rect 379 94 387 99
rect 379 92 382 94
rect 384 92 387 94
rect 379 90 387 92
rect 389 94 396 103
rect 389 92 392 94
rect 394 92 396 94
rect 389 90 396 92
rect 411 83 416 104
rect 418 94 432 110
rect 418 92 421 94
rect 423 92 432 94
rect 434 108 442 110
rect 434 106 437 108
rect 439 106 442 108
rect 434 101 442 106
rect 434 99 437 101
rect 439 99 442 101
rect 434 92 442 99
rect 444 101 452 110
rect 444 99 447 101
rect 449 99 452 101
rect 444 92 452 99
rect 418 87 430 92
rect 418 85 421 87
rect 423 85 430 87
rect 418 83 430 85
rect 447 83 452 92
rect 454 95 459 110
rect 467 106 472 111
rect 465 104 472 106
rect 465 102 467 104
rect 469 102 472 104
rect 465 97 472 102
rect 465 95 467 97
rect 469 95 472 97
rect 454 93 461 95
rect 465 93 472 95
rect 474 104 482 111
rect 505 108 512 110
rect 505 106 507 108
rect 509 106 512 108
rect 474 93 485 104
rect 454 91 457 93
rect 459 91 461 93
rect 454 89 461 91
rect 454 83 459 89
rect 476 87 485 93
rect 476 85 478 87
rect 480 85 485 87
rect 476 83 485 85
rect 487 83 492 104
rect 494 96 499 104
rect 505 101 512 106
rect 505 99 507 101
rect 509 99 512 101
rect 505 97 512 99
rect 494 94 501 96
rect 494 92 497 94
rect 499 92 501 94
rect 507 92 512 97
rect 514 103 520 110
rect 554 108 561 110
rect 554 106 556 108
rect 558 106 561 108
rect 554 104 561 106
rect 514 96 522 103
rect 514 94 517 96
rect 519 94 522 96
rect 514 92 522 94
rect 494 90 501 92
rect 494 83 499 90
rect 516 90 522 92
rect 524 101 532 103
rect 524 99 527 101
rect 529 99 532 101
rect 524 94 532 99
rect 524 92 527 94
rect 529 92 532 94
rect 524 90 532 92
rect 534 94 541 103
rect 534 92 537 94
rect 539 92 541 94
rect 534 90 541 92
rect 556 83 561 104
rect 563 94 577 110
rect 563 92 566 94
rect 568 92 577 94
rect 579 108 587 110
rect 579 106 582 108
rect 584 106 587 108
rect 579 101 587 106
rect 579 99 582 101
rect 584 99 587 101
rect 579 92 587 99
rect 589 101 597 110
rect 589 99 592 101
rect 594 99 597 101
rect 589 92 597 99
rect 563 87 575 92
rect 563 85 566 87
rect 568 85 575 87
rect 563 83 575 85
rect 592 83 597 92
rect 599 95 604 110
rect 610 108 617 110
rect 610 106 612 108
rect 614 106 617 108
rect 610 101 617 106
rect 610 99 612 101
rect 614 99 617 101
rect 610 97 617 99
rect 599 93 606 95
rect 599 91 602 93
rect 604 91 606 93
rect 612 92 617 97
rect 619 103 625 110
rect 659 108 666 110
rect 659 106 661 108
rect 663 106 666 108
rect 659 104 666 106
rect 619 96 627 103
rect 619 94 622 96
rect 624 94 627 96
rect 619 92 627 94
rect 599 89 606 91
rect 599 83 604 89
rect 621 90 627 92
rect 629 101 637 103
rect 629 99 632 101
rect 634 99 637 101
rect 629 94 637 99
rect 629 92 632 94
rect 634 92 637 94
rect 629 90 637 92
rect 639 94 646 103
rect 639 92 642 94
rect 644 92 646 94
rect 639 90 646 92
rect 661 83 666 104
rect 668 94 682 110
rect 668 92 671 94
rect 673 92 682 94
rect 684 108 692 110
rect 684 106 687 108
rect 689 106 692 108
rect 684 101 692 106
rect 684 99 687 101
rect 689 99 692 101
rect 684 92 692 99
rect 694 101 702 110
rect 694 99 697 101
rect 699 99 702 101
rect 694 92 702 99
rect 668 87 680 92
rect 668 85 671 87
rect 673 85 680 87
rect 668 83 680 85
rect 697 83 702 92
rect 704 95 709 110
rect 717 106 722 111
rect 715 104 722 106
rect 715 102 717 104
rect 719 102 722 104
rect 715 97 722 102
rect 715 95 717 97
rect 719 95 722 97
rect 704 93 711 95
rect 715 93 722 95
rect 724 104 732 111
rect 755 108 762 110
rect 755 106 757 108
rect 759 106 762 108
rect 724 93 735 104
rect 704 91 707 93
rect 709 91 711 93
rect 704 89 711 91
rect 704 83 709 89
rect 726 87 735 93
rect 726 85 728 87
rect 730 85 735 87
rect 726 83 735 85
rect 737 83 742 104
rect 744 96 749 104
rect 755 101 762 106
rect 755 99 757 101
rect 759 99 762 101
rect 755 97 762 99
rect 744 94 751 96
rect 744 92 747 94
rect 749 92 751 94
rect 757 92 762 97
rect 764 103 770 110
rect 804 108 811 110
rect 804 106 806 108
rect 808 106 811 108
rect 804 104 811 106
rect 764 96 772 103
rect 764 94 767 96
rect 769 94 772 96
rect 764 92 772 94
rect 744 90 751 92
rect 744 83 749 90
rect 766 90 772 92
rect 774 101 782 103
rect 774 99 777 101
rect 779 99 782 101
rect 774 94 782 99
rect 774 92 777 94
rect 779 92 782 94
rect 774 90 782 92
rect 784 94 791 103
rect 784 92 787 94
rect 789 92 791 94
rect 784 90 791 92
rect 806 83 811 104
rect 813 94 827 110
rect 813 92 816 94
rect 818 92 827 94
rect 829 108 837 110
rect 829 106 832 108
rect 834 106 837 108
rect 829 101 837 106
rect 829 99 832 101
rect 834 99 837 101
rect 829 92 837 99
rect 839 101 847 110
rect 839 99 842 101
rect 844 99 847 101
rect 839 92 847 99
rect 813 87 825 92
rect 813 85 816 87
rect 818 85 825 87
rect 813 83 825 85
rect 842 83 847 92
rect 849 95 854 110
rect 860 108 867 110
rect 860 106 862 108
rect 864 106 867 108
rect 860 101 867 106
rect 860 99 862 101
rect 864 99 867 101
rect 860 97 867 99
rect 849 93 856 95
rect 849 91 852 93
rect 854 91 856 93
rect 862 92 867 97
rect 869 103 875 110
rect 909 108 916 110
rect 909 106 911 108
rect 913 106 916 108
rect 909 104 916 106
rect 869 96 877 103
rect 869 94 872 96
rect 874 94 877 96
rect 869 92 877 94
rect 849 89 856 91
rect 849 83 854 89
rect 871 90 877 92
rect 879 101 887 103
rect 879 99 882 101
rect 884 99 887 101
rect 879 94 887 99
rect 879 92 882 94
rect 884 92 887 94
rect 879 90 887 92
rect 889 94 896 103
rect 889 92 892 94
rect 894 92 896 94
rect 889 90 896 92
rect 911 83 916 104
rect 918 94 932 110
rect 918 92 921 94
rect 923 92 932 94
rect 934 108 942 110
rect 934 106 937 108
rect 939 106 942 108
rect 934 101 942 106
rect 934 99 937 101
rect 939 99 942 101
rect 934 92 942 99
rect 944 101 952 110
rect 944 99 947 101
rect 949 99 952 101
rect 944 92 952 99
rect 918 87 930 92
rect 918 85 921 87
rect 923 85 930 87
rect 918 83 930 85
rect 947 83 952 92
rect 954 95 959 110
rect 967 106 972 111
rect 965 104 972 106
rect 965 102 967 104
rect 969 102 972 104
rect 965 97 972 102
rect 965 95 967 97
rect 969 95 972 97
rect 954 93 961 95
rect 965 93 972 95
rect 974 104 982 111
rect 1005 108 1012 110
rect 1005 106 1007 108
rect 1009 106 1012 108
rect 974 93 985 104
rect 954 91 957 93
rect 959 91 961 93
rect 954 89 961 91
rect 954 83 959 89
rect 976 87 985 93
rect 976 85 978 87
rect 980 85 985 87
rect 976 83 985 85
rect 987 83 992 104
rect 994 96 999 104
rect 1005 101 1012 106
rect 1005 99 1007 101
rect 1009 99 1012 101
rect 1005 97 1012 99
rect 994 94 1001 96
rect 994 92 997 94
rect 999 92 1001 94
rect 1007 92 1012 97
rect 1014 103 1020 110
rect 1054 108 1061 110
rect 1054 106 1056 108
rect 1058 106 1061 108
rect 1054 104 1061 106
rect 1014 96 1022 103
rect 1014 94 1017 96
rect 1019 94 1022 96
rect 1014 92 1022 94
rect 994 90 1001 92
rect 994 83 999 90
rect 1016 90 1022 92
rect 1024 101 1032 103
rect 1024 99 1027 101
rect 1029 99 1032 101
rect 1024 94 1032 99
rect 1024 92 1027 94
rect 1029 92 1032 94
rect 1024 90 1032 92
rect 1034 94 1041 103
rect 1034 92 1037 94
rect 1039 92 1041 94
rect 1034 90 1041 92
rect 1056 83 1061 104
rect 1063 94 1077 110
rect 1063 92 1066 94
rect 1068 92 1077 94
rect 1079 108 1087 110
rect 1079 106 1082 108
rect 1084 106 1087 108
rect 1079 101 1087 106
rect 1079 99 1082 101
rect 1084 99 1087 101
rect 1079 92 1087 99
rect 1089 101 1097 110
rect 1089 99 1092 101
rect 1094 99 1097 101
rect 1089 92 1097 99
rect 1063 87 1075 92
rect 1063 85 1066 87
rect 1068 85 1075 87
rect 1063 83 1075 85
rect 1092 83 1097 92
rect 1099 95 1104 110
rect 1110 108 1117 110
rect 1110 106 1112 108
rect 1114 106 1117 108
rect 1110 101 1117 106
rect 1110 99 1112 101
rect 1114 99 1117 101
rect 1110 97 1117 99
rect 1099 93 1106 95
rect 1099 91 1102 93
rect 1104 91 1106 93
rect 1112 92 1117 97
rect 1119 103 1125 110
rect 1159 108 1166 110
rect 1159 106 1161 108
rect 1163 106 1166 108
rect 1159 104 1166 106
rect 1119 96 1127 103
rect 1119 94 1122 96
rect 1124 94 1127 96
rect 1119 92 1127 94
rect 1099 89 1106 91
rect 1099 83 1104 89
rect 1121 90 1127 92
rect 1129 101 1137 103
rect 1129 99 1132 101
rect 1134 99 1137 101
rect 1129 94 1137 99
rect 1129 92 1132 94
rect 1134 92 1137 94
rect 1129 90 1137 92
rect 1139 94 1146 103
rect 1139 92 1142 94
rect 1144 92 1146 94
rect 1139 90 1146 92
rect 1161 83 1166 104
rect 1168 94 1182 110
rect 1168 92 1171 94
rect 1173 92 1182 94
rect 1184 108 1192 110
rect 1184 106 1187 108
rect 1189 106 1192 108
rect 1184 101 1192 106
rect 1184 99 1187 101
rect 1189 99 1192 101
rect 1184 92 1192 99
rect 1194 101 1202 110
rect 1194 99 1197 101
rect 1199 99 1202 101
rect 1194 92 1202 99
rect 1168 87 1180 92
rect 1168 85 1171 87
rect 1173 85 1180 87
rect 1168 83 1180 85
rect 1197 83 1202 92
rect 1204 95 1209 110
rect 1204 93 1211 95
rect 1204 91 1207 93
rect 1209 91 1211 93
rect 1204 89 1211 91
rect 1204 83 1209 89
rect 18 69 27 71
rect 18 67 20 69
rect 22 67 27 69
rect 18 61 27 67
rect 7 59 14 61
rect 7 57 9 59
rect 11 57 14 59
rect 7 52 14 57
rect 7 50 9 52
rect 11 50 14 52
rect 7 48 14 50
rect 9 43 14 48
rect 16 50 27 61
rect 29 50 34 71
rect 36 64 41 71
rect 36 62 43 64
rect 58 62 64 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 58 43 60
rect 36 50 41 58
rect 49 57 54 62
rect 47 55 54 57
rect 47 53 49 55
rect 51 53 54 55
rect 16 43 24 50
rect 47 48 54 53
rect 47 46 49 48
rect 51 46 54 48
rect 47 44 54 46
rect 56 60 64 62
rect 56 58 59 60
rect 61 58 64 60
rect 56 51 64 58
rect 66 62 74 64
rect 66 60 69 62
rect 71 60 74 62
rect 66 55 74 60
rect 66 53 69 55
rect 71 53 74 55
rect 66 51 74 53
rect 76 62 83 64
rect 76 60 79 62
rect 81 60 83 62
rect 76 51 83 60
rect 56 44 62 51
rect 98 50 103 71
rect 96 48 103 50
rect 96 46 98 48
rect 100 46 103 48
rect 96 44 103 46
rect 105 69 117 71
rect 105 67 108 69
rect 110 67 117 69
rect 105 62 117 67
rect 134 62 139 71
rect 105 60 108 62
rect 110 60 119 62
rect 105 44 119 60
rect 121 55 129 62
rect 121 53 124 55
rect 126 53 129 55
rect 121 48 129 53
rect 121 46 124 48
rect 126 46 129 48
rect 121 44 129 46
rect 131 55 139 62
rect 131 53 134 55
rect 136 53 139 55
rect 131 44 139 53
rect 141 65 146 71
rect 141 63 148 65
rect 141 61 144 63
rect 146 61 148 63
rect 163 62 169 64
rect 141 59 148 61
rect 141 44 146 59
rect 154 57 159 62
rect 152 55 159 57
rect 152 53 154 55
rect 156 53 159 55
rect 152 48 159 53
rect 152 46 154 48
rect 156 46 159 48
rect 152 44 159 46
rect 161 60 169 62
rect 161 58 164 60
rect 166 58 169 60
rect 161 51 169 58
rect 171 62 179 64
rect 171 60 174 62
rect 176 60 179 62
rect 171 55 179 60
rect 171 53 174 55
rect 176 53 179 55
rect 171 51 179 53
rect 181 62 188 64
rect 181 60 184 62
rect 186 60 188 62
rect 181 51 188 60
rect 161 44 167 51
rect 203 50 208 71
rect 201 48 208 50
rect 201 46 203 48
rect 205 46 208 48
rect 201 44 208 46
rect 210 69 222 71
rect 210 67 213 69
rect 215 67 222 69
rect 210 62 222 67
rect 239 62 244 71
rect 210 60 213 62
rect 215 60 224 62
rect 210 44 224 60
rect 226 55 234 62
rect 226 53 229 55
rect 231 53 234 55
rect 226 48 234 53
rect 226 46 229 48
rect 231 46 234 48
rect 226 44 234 46
rect 236 55 244 62
rect 236 53 239 55
rect 241 53 244 55
rect 236 44 244 53
rect 246 65 251 71
rect 268 69 277 71
rect 268 67 270 69
rect 272 67 277 69
rect 246 63 253 65
rect 246 61 249 63
rect 251 61 253 63
rect 268 61 277 67
rect 246 59 253 61
rect 257 59 264 61
rect 246 44 251 59
rect 257 57 259 59
rect 261 57 264 59
rect 257 52 264 57
rect 257 50 259 52
rect 261 50 264 52
rect 257 48 264 50
rect 259 43 264 48
rect 266 50 277 61
rect 279 50 284 71
rect 286 64 291 71
rect 286 62 293 64
rect 308 62 314 64
rect 286 60 289 62
rect 291 60 293 62
rect 286 58 293 60
rect 286 50 291 58
rect 299 57 304 62
rect 297 55 304 57
rect 297 53 299 55
rect 301 53 304 55
rect 266 43 274 50
rect 297 48 304 53
rect 297 46 299 48
rect 301 46 304 48
rect 297 44 304 46
rect 306 60 314 62
rect 306 58 309 60
rect 311 58 314 60
rect 306 51 314 58
rect 316 62 324 64
rect 316 60 319 62
rect 321 60 324 62
rect 316 55 324 60
rect 316 53 319 55
rect 321 53 324 55
rect 316 51 324 53
rect 326 62 333 64
rect 326 60 329 62
rect 331 60 333 62
rect 326 51 333 60
rect 306 44 312 51
rect 348 50 353 71
rect 346 48 353 50
rect 346 46 348 48
rect 350 46 353 48
rect 346 44 353 46
rect 355 69 367 71
rect 355 67 358 69
rect 360 67 367 69
rect 355 62 367 67
rect 384 62 389 71
rect 355 60 358 62
rect 360 60 369 62
rect 355 44 369 60
rect 371 55 379 62
rect 371 53 374 55
rect 376 53 379 55
rect 371 48 379 53
rect 371 46 374 48
rect 376 46 379 48
rect 371 44 379 46
rect 381 55 389 62
rect 381 53 384 55
rect 386 53 389 55
rect 381 44 389 53
rect 391 65 396 71
rect 391 63 398 65
rect 391 61 394 63
rect 396 61 398 63
rect 413 62 419 64
rect 391 59 398 61
rect 391 44 396 59
rect 404 57 409 62
rect 402 55 409 57
rect 402 53 404 55
rect 406 53 409 55
rect 402 48 409 53
rect 402 46 404 48
rect 406 46 409 48
rect 402 44 409 46
rect 411 60 419 62
rect 411 58 414 60
rect 416 58 419 60
rect 411 51 419 58
rect 421 62 429 64
rect 421 60 424 62
rect 426 60 429 62
rect 421 55 429 60
rect 421 53 424 55
rect 426 53 429 55
rect 421 51 429 53
rect 431 62 438 64
rect 431 60 434 62
rect 436 60 438 62
rect 431 51 438 60
rect 411 44 417 51
rect 453 50 458 71
rect 451 48 458 50
rect 451 46 453 48
rect 455 46 458 48
rect 451 44 458 46
rect 460 69 472 71
rect 460 67 463 69
rect 465 67 472 69
rect 460 62 472 67
rect 489 62 494 71
rect 460 60 463 62
rect 465 60 474 62
rect 460 44 474 60
rect 476 55 484 62
rect 476 53 479 55
rect 481 53 484 55
rect 476 48 484 53
rect 476 46 479 48
rect 481 46 484 48
rect 476 44 484 46
rect 486 55 494 62
rect 486 53 489 55
rect 491 53 494 55
rect 486 44 494 53
rect 496 65 501 71
rect 518 69 527 71
rect 518 67 520 69
rect 522 67 527 69
rect 496 63 503 65
rect 496 61 499 63
rect 501 61 503 63
rect 518 61 527 67
rect 496 59 503 61
rect 507 59 514 61
rect 496 44 501 59
rect 507 57 509 59
rect 511 57 514 59
rect 507 52 514 57
rect 507 50 509 52
rect 511 50 514 52
rect 507 48 514 50
rect 509 43 514 48
rect 516 50 527 61
rect 529 50 534 71
rect 536 64 541 71
rect 536 62 543 64
rect 558 62 564 64
rect 536 60 539 62
rect 541 60 543 62
rect 536 58 543 60
rect 536 50 541 58
rect 549 57 554 62
rect 547 55 554 57
rect 547 53 549 55
rect 551 53 554 55
rect 516 43 524 50
rect 547 48 554 53
rect 547 46 549 48
rect 551 46 554 48
rect 547 44 554 46
rect 556 60 564 62
rect 556 58 559 60
rect 561 58 564 60
rect 556 51 564 58
rect 566 62 574 64
rect 566 60 569 62
rect 571 60 574 62
rect 566 55 574 60
rect 566 53 569 55
rect 571 53 574 55
rect 566 51 574 53
rect 576 62 583 64
rect 576 60 579 62
rect 581 60 583 62
rect 576 51 583 60
rect 556 44 562 51
rect 598 50 603 71
rect 596 48 603 50
rect 596 46 598 48
rect 600 46 603 48
rect 596 44 603 46
rect 605 69 617 71
rect 605 67 608 69
rect 610 67 617 69
rect 605 62 617 67
rect 634 62 639 71
rect 605 60 608 62
rect 610 60 619 62
rect 605 44 619 60
rect 621 55 629 62
rect 621 53 624 55
rect 626 53 629 55
rect 621 48 629 53
rect 621 46 624 48
rect 626 46 629 48
rect 621 44 629 46
rect 631 55 639 62
rect 631 53 634 55
rect 636 53 639 55
rect 631 44 639 53
rect 641 65 646 71
rect 641 63 648 65
rect 641 61 644 63
rect 646 61 648 63
rect 663 62 669 64
rect 641 59 648 61
rect 641 44 646 59
rect 654 57 659 62
rect 652 55 659 57
rect 652 53 654 55
rect 656 53 659 55
rect 652 48 659 53
rect 652 46 654 48
rect 656 46 659 48
rect 652 44 659 46
rect 661 60 669 62
rect 661 58 664 60
rect 666 58 669 60
rect 661 51 669 58
rect 671 62 679 64
rect 671 60 674 62
rect 676 60 679 62
rect 671 55 679 60
rect 671 53 674 55
rect 676 53 679 55
rect 671 51 679 53
rect 681 62 688 64
rect 681 60 684 62
rect 686 60 688 62
rect 681 51 688 60
rect 661 44 667 51
rect 703 50 708 71
rect 701 48 708 50
rect 701 46 703 48
rect 705 46 708 48
rect 701 44 708 46
rect 710 69 722 71
rect 710 67 713 69
rect 715 67 722 69
rect 710 62 722 67
rect 739 62 744 71
rect 710 60 713 62
rect 715 60 724 62
rect 710 44 724 60
rect 726 55 734 62
rect 726 53 729 55
rect 731 53 734 55
rect 726 48 734 53
rect 726 46 729 48
rect 731 46 734 48
rect 726 44 734 46
rect 736 55 744 62
rect 736 53 739 55
rect 741 53 744 55
rect 736 44 744 53
rect 746 65 751 71
rect 768 69 777 71
rect 768 67 770 69
rect 772 67 777 69
rect 746 63 753 65
rect 746 61 749 63
rect 751 61 753 63
rect 768 61 777 67
rect 746 59 753 61
rect 757 59 764 61
rect 746 44 751 59
rect 757 57 759 59
rect 761 57 764 59
rect 757 52 764 57
rect 757 50 759 52
rect 761 50 764 52
rect 757 48 764 50
rect 759 43 764 48
rect 766 50 777 61
rect 779 50 784 71
rect 786 64 791 71
rect 786 62 793 64
rect 808 62 814 64
rect 786 60 789 62
rect 791 60 793 62
rect 786 58 793 60
rect 786 50 791 58
rect 799 57 804 62
rect 797 55 804 57
rect 797 53 799 55
rect 801 53 804 55
rect 766 43 774 50
rect 797 48 804 53
rect 797 46 799 48
rect 801 46 804 48
rect 797 44 804 46
rect 806 60 814 62
rect 806 58 809 60
rect 811 58 814 60
rect 806 51 814 58
rect 816 62 824 64
rect 816 60 819 62
rect 821 60 824 62
rect 816 55 824 60
rect 816 53 819 55
rect 821 53 824 55
rect 816 51 824 53
rect 826 62 833 64
rect 826 60 829 62
rect 831 60 833 62
rect 826 51 833 60
rect 806 44 812 51
rect 848 50 853 71
rect 846 48 853 50
rect 846 46 848 48
rect 850 46 853 48
rect 846 44 853 46
rect 855 69 867 71
rect 855 67 858 69
rect 860 67 867 69
rect 855 62 867 67
rect 884 62 889 71
rect 855 60 858 62
rect 860 60 869 62
rect 855 44 869 60
rect 871 55 879 62
rect 871 53 874 55
rect 876 53 879 55
rect 871 48 879 53
rect 871 46 874 48
rect 876 46 879 48
rect 871 44 879 46
rect 881 55 889 62
rect 881 53 884 55
rect 886 53 889 55
rect 881 44 889 53
rect 891 65 896 71
rect 891 63 898 65
rect 891 61 894 63
rect 896 61 898 63
rect 913 62 919 64
rect 891 59 898 61
rect 891 44 896 59
rect 904 57 909 62
rect 902 55 909 57
rect 902 53 904 55
rect 906 53 909 55
rect 902 48 909 53
rect 902 46 904 48
rect 906 46 909 48
rect 902 44 909 46
rect 911 60 919 62
rect 911 58 914 60
rect 916 58 919 60
rect 911 51 919 58
rect 921 62 929 64
rect 921 60 924 62
rect 926 60 929 62
rect 921 55 929 60
rect 921 53 924 55
rect 926 53 929 55
rect 921 51 929 53
rect 931 62 938 64
rect 931 60 934 62
rect 936 60 938 62
rect 931 51 938 60
rect 911 44 917 51
rect 953 50 958 71
rect 951 48 958 50
rect 951 46 953 48
rect 955 46 958 48
rect 951 44 958 46
rect 960 69 972 71
rect 960 67 963 69
rect 965 67 972 69
rect 960 62 972 67
rect 989 62 994 71
rect 960 60 963 62
rect 965 60 974 62
rect 960 44 974 60
rect 976 55 984 62
rect 976 53 979 55
rect 981 53 984 55
rect 976 48 984 53
rect 976 46 979 48
rect 981 46 984 48
rect 976 44 984 46
rect 986 55 994 62
rect 986 53 989 55
rect 991 53 994 55
rect 986 44 994 53
rect 996 65 1001 71
rect 996 63 1003 65
rect 996 61 999 63
rect 1001 61 1003 63
rect 996 59 1003 61
rect 996 44 1001 59
<< alu1 >>
rect 4 413 202 418
rect 4 411 35 413
rect 37 411 45 413
rect 47 411 75 413
rect 77 411 85 413
rect 87 411 103 413
rect 105 411 156 413
rect 158 411 187 413
rect 189 411 197 413
rect 199 411 202 413
rect 486 415 889 420
rect 486 413 517 415
rect 519 413 527 415
rect 529 413 557 415
rect 559 413 567 415
rect 569 413 585 415
rect 587 413 638 415
rect 640 413 669 415
rect 671 413 679 415
rect 681 413 722 415
rect 724 413 732 415
rect 734 413 762 415
rect 764 413 772 415
rect 774 413 790 415
rect 792 413 843 415
rect 845 413 874 415
rect 876 413 884 415
rect 886 413 889 415
rect 486 412 889 413
rect 4 410 202 411
rect 21 388 26 397
rect 38 401 50 405
rect 38 399 46 401
rect 48 399 50 401
rect 46 396 50 399
rect 21 387 35 388
rect 21 385 29 387
rect 31 385 32 387
rect 34 385 35 387
rect 21 384 35 385
rect 14 379 27 380
rect 14 377 19 379
rect 21 377 27 379
rect 14 376 27 377
rect 14 371 18 376
rect 46 394 47 396
rect 49 394 50 396
rect 46 379 50 394
rect 61 388 66 397
rect 78 401 90 405
rect 78 399 86 401
rect 88 399 90 401
rect 61 387 75 388
rect 61 385 69 387
rect 71 385 72 387
rect 74 385 75 387
rect 61 384 75 385
rect 14 369 15 371
rect 17 369 18 371
rect 14 367 18 369
rect 45 377 50 379
rect 45 375 46 377
rect 48 375 50 377
rect 45 370 50 375
rect 45 368 46 370
rect 48 368 50 370
rect 45 366 50 368
rect 54 379 67 380
rect 54 377 59 379
rect 61 377 67 379
rect 54 376 67 377
rect 54 372 58 376
rect 86 379 90 399
rect 54 370 55 372
rect 57 370 58 372
rect 54 367 58 370
rect 85 377 90 379
rect 85 375 86 377
rect 88 375 90 377
rect 85 373 90 375
rect 85 371 86 373
rect 88 371 90 373
rect 85 370 90 371
rect 85 368 86 370
rect 88 368 90 370
rect 85 366 90 368
rect 101 403 125 404
rect 101 401 121 403
rect 123 401 125 403
rect 101 400 125 401
rect 101 372 105 400
rect 140 396 153 397
rect 140 394 148 396
rect 150 394 153 396
rect 140 392 153 394
rect 140 390 141 392
rect 143 391 153 392
rect 143 390 145 391
rect 101 370 117 372
rect 101 368 113 370
rect 115 368 117 370
rect 101 367 117 368
rect 140 383 145 390
rect 173 396 178 397
rect 173 394 175 396
rect 177 394 178 396
rect 173 388 178 394
rect 190 401 202 405
rect 190 399 198 401
rect 200 399 202 401
rect 173 387 187 388
rect 173 385 181 387
rect 183 385 187 387
rect 173 384 187 385
rect 156 380 161 381
rect 156 379 162 380
rect 166 379 179 380
rect 156 377 157 379
rect 159 377 171 379
rect 173 377 179 379
rect 156 376 179 377
rect 156 374 170 376
rect 156 365 161 374
rect 166 373 170 374
rect 198 384 202 399
rect 503 390 508 399
rect 520 403 532 407
rect 520 401 528 403
rect 530 401 532 403
rect 528 398 532 401
rect 503 389 517 390
rect 503 387 511 389
rect 513 387 514 389
rect 516 387 517 389
rect 503 386 517 387
rect 198 382 199 384
rect 201 382 202 384
rect 198 379 202 382
rect 166 371 167 373
rect 169 371 170 373
rect 166 367 170 371
rect 197 377 202 379
rect 197 375 198 377
rect 200 375 202 377
rect 197 370 202 375
rect 149 359 161 365
rect 197 368 198 370
rect 200 368 202 370
rect 496 381 509 382
rect 496 379 501 381
rect 503 379 509 381
rect 496 378 509 379
rect 496 373 500 378
rect 528 396 529 398
rect 531 396 532 398
rect 528 381 532 396
rect 543 390 548 399
rect 560 403 572 407
rect 560 401 568 403
rect 570 401 572 403
rect 543 389 557 390
rect 543 387 551 389
rect 553 387 554 389
rect 556 387 557 389
rect 543 386 557 387
rect 496 371 497 373
rect 499 371 500 373
rect 496 369 500 371
rect 527 379 532 381
rect 527 377 528 379
rect 530 377 532 379
rect 527 372 532 377
rect 197 366 202 368
rect 527 370 528 372
rect 530 370 532 372
rect 527 368 532 370
rect 536 381 549 382
rect 536 379 541 381
rect 543 379 549 381
rect 536 378 549 379
rect 536 374 540 378
rect 568 381 572 401
rect 536 372 537 374
rect 539 372 540 374
rect 536 369 540 372
rect 567 379 572 381
rect 567 377 568 379
rect 570 377 572 379
rect 567 375 572 377
rect 567 373 568 375
rect 570 373 572 375
rect 567 372 572 373
rect 567 370 568 372
rect 570 370 572 372
rect 567 368 572 370
rect 583 405 607 406
rect 583 403 603 405
rect 605 403 607 405
rect 583 402 607 403
rect 583 374 587 402
rect 622 398 635 399
rect 622 396 630 398
rect 632 396 635 398
rect 622 394 635 396
rect 622 392 623 394
rect 625 393 635 394
rect 625 392 627 393
rect 583 372 599 374
rect 583 370 595 372
rect 597 370 599 372
rect 583 369 599 370
rect 622 385 627 392
rect 655 398 660 399
rect 655 396 657 398
rect 659 396 660 398
rect 655 390 660 396
rect 672 403 684 407
rect 672 401 680 403
rect 682 401 684 403
rect 655 389 669 390
rect 655 387 663 389
rect 665 387 669 389
rect 655 386 669 387
rect 638 382 643 383
rect 638 381 644 382
rect 648 381 661 382
rect 638 379 639 381
rect 641 379 653 381
rect 655 379 661 381
rect 638 378 661 379
rect 638 376 652 378
rect 638 367 643 376
rect 648 375 652 376
rect 680 386 684 401
rect 708 390 713 399
rect 725 403 737 407
rect 725 401 733 403
rect 735 401 737 403
rect 733 398 737 401
rect 708 389 722 390
rect 708 387 716 389
rect 718 387 719 389
rect 721 387 722 389
rect 708 386 722 387
rect 680 384 681 386
rect 683 384 684 386
rect 680 381 684 384
rect 648 373 649 375
rect 651 373 652 375
rect 648 369 652 373
rect 679 379 684 381
rect 679 377 680 379
rect 682 377 684 379
rect 679 372 684 377
rect 631 361 643 367
rect 679 370 680 372
rect 682 370 684 372
rect 679 368 684 370
rect 701 381 714 382
rect 701 379 706 381
rect 708 379 714 381
rect 701 378 714 379
rect 701 373 705 378
rect 733 396 734 398
rect 736 396 737 398
rect 733 381 737 396
rect 748 390 753 399
rect 765 403 777 407
rect 765 401 773 403
rect 775 401 777 403
rect 748 389 762 390
rect 748 387 756 389
rect 758 387 759 389
rect 761 387 762 389
rect 748 386 762 387
rect 701 371 702 373
rect 704 371 705 373
rect 701 369 705 371
rect 732 379 737 381
rect 732 377 733 379
rect 735 377 737 379
rect 732 372 737 377
rect 732 370 733 372
rect 735 370 737 372
rect 732 368 737 370
rect 741 381 754 382
rect 741 379 746 381
rect 748 379 754 381
rect 741 378 754 379
rect 741 374 745 378
rect 773 381 777 401
rect 741 372 742 374
rect 744 372 745 374
rect 741 369 745 372
rect 772 379 777 381
rect 772 377 773 379
rect 775 377 777 379
rect 772 375 777 377
rect 772 373 773 375
rect 775 373 777 375
rect 772 372 777 373
rect 772 370 773 372
rect 775 370 777 372
rect 772 368 777 370
rect 788 405 812 406
rect 788 403 808 405
rect 810 403 812 405
rect 788 402 812 403
rect 788 374 792 402
rect 827 398 840 399
rect 827 396 835 398
rect 837 396 840 398
rect 827 394 840 396
rect 827 392 828 394
rect 830 393 840 394
rect 830 392 832 393
rect 788 372 804 374
rect 788 370 800 372
rect 802 370 804 372
rect 788 369 804 370
rect 827 385 832 392
rect 860 398 865 399
rect 860 396 862 398
rect 864 396 865 398
rect 860 390 865 396
rect 877 403 889 407
rect 877 401 885 403
rect 887 401 889 403
rect 860 389 874 390
rect 860 387 868 389
rect 870 387 874 389
rect 860 386 874 387
rect 843 382 848 383
rect 843 381 849 382
rect 853 381 866 382
rect 843 379 844 381
rect 846 379 858 381
rect 860 379 866 381
rect 843 378 866 379
rect 843 376 857 378
rect 843 367 848 376
rect 853 375 857 376
rect 885 386 889 401
rect 885 384 886 386
rect 888 384 889 386
rect 885 381 889 384
rect 853 373 854 375
rect 856 373 857 375
rect 853 369 857 373
rect 884 379 889 381
rect 884 377 885 379
rect 887 377 889 379
rect 884 372 889 377
rect 836 361 848 367
rect 884 370 885 372
rect 887 370 889 372
rect 884 368 889 370
rect 495 355 889 356
rect 13 353 202 354
rect 13 351 45 353
rect 47 351 85 353
rect 87 351 123 353
rect 125 351 197 353
rect 199 351 202 353
rect 13 341 202 351
rect 13 339 17 341
rect 19 339 85 341
rect 87 339 97 341
rect 99 339 171 341
rect 173 339 202 341
rect 495 353 527 355
rect 529 353 567 355
rect 569 353 605 355
rect 607 353 679 355
rect 681 353 732 355
rect 734 353 772 355
rect 774 353 810 355
rect 812 353 884 355
rect 886 353 889 355
rect 495 343 889 353
rect 495 341 499 343
rect 501 341 567 343
rect 569 341 579 343
rect 581 341 653 343
rect 655 341 704 343
rect 706 341 772 343
rect 774 341 784 343
rect 786 341 858 343
rect 860 341 889 343
rect 495 340 889 341
rect 13 338 202 339
rect 14 324 19 326
rect 14 322 16 324
rect 18 322 19 324
rect 14 317 19 322
rect 14 315 16 317
rect 18 315 19 317
rect 14 313 19 315
rect 46 324 50 325
rect 46 322 47 324
rect 49 322 50 324
rect 14 293 18 313
rect 46 316 50 322
rect 37 315 50 316
rect 37 313 43 315
rect 45 313 50 315
rect 37 312 50 313
rect 54 316 58 325
rect 85 324 90 326
rect 54 315 67 316
rect 54 313 55 315
rect 57 313 59 315
rect 61 313 67 315
rect 54 312 67 313
rect 29 307 43 308
rect 29 305 30 307
rect 32 305 33 307
rect 35 305 43 307
rect 29 304 43 305
rect 14 291 16 293
rect 18 291 26 293
rect 14 287 26 291
rect 38 295 43 304
rect 61 307 75 308
rect 61 305 69 307
rect 71 305 72 307
rect 74 305 75 307
rect 61 304 75 305
rect 85 322 86 324
rect 88 322 90 324
rect 85 317 90 322
rect 85 315 86 317
rect 88 315 90 317
rect 85 313 90 315
rect 61 295 66 304
rect 86 298 90 313
rect 86 296 87 298
rect 89 296 90 298
rect 86 293 90 296
rect 78 291 86 293
rect 88 291 90 293
rect 78 287 90 291
rect 94 324 99 326
rect 94 322 96 324
rect 98 322 99 324
rect 135 331 147 333
rect 135 329 143 331
rect 145 329 147 331
rect 135 327 147 329
rect 94 317 99 322
rect 94 315 96 317
rect 98 315 99 317
rect 94 313 99 315
rect 94 293 98 313
rect 126 318 130 325
rect 135 318 140 327
rect 496 326 501 328
rect 126 316 140 318
rect 117 315 140 316
rect 117 313 123 315
rect 125 313 137 315
rect 139 313 140 315
rect 117 312 130 313
rect 134 312 140 313
rect 135 311 140 312
rect 109 307 123 308
rect 109 305 113 307
rect 115 305 123 307
rect 109 304 123 305
rect 94 291 96 293
rect 98 291 106 293
rect 94 287 106 291
rect 118 298 123 304
rect 118 296 119 298
rect 121 296 123 298
rect 118 295 123 296
rect 151 302 156 309
rect 179 324 195 325
rect 179 322 181 324
rect 183 322 195 324
rect 179 320 195 322
rect 151 301 153 302
rect 143 300 153 301
rect 155 300 156 302
rect 143 298 156 300
rect 143 296 146 298
rect 148 296 156 298
rect 143 295 156 296
rect 191 292 195 320
rect 171 291 195 292
rect 171 289 173 291
rect 175 289 195 291
rect 496 324 498 326
rect 500 324 501 326
rect 496 319 501 324
rect 496 317 498 319
rect 500 317 501 319
rect 496 315 501 317
rect 528 326 532 327
rect 528 324 529 326
rect 531 324 532 326
rect 496 295 500 315
rect 528 318 532 324
rect 519 317 532 318
rect 519 315 525 317
rect 527 315 532 317
rect 519 314 532 315
rect 536 318 540 327
rect 567 326 572 328
rect 536 317 549 318
rect 536 315 537 317
rect 539 315 541 317
rect 543 315 549 317
rect 536 314 549 315
rect 511 309 525 310
rect 511 307 512 309
rect 514 307 515 309
rect 517 307 525 309
rect 511 306 525 307
rect 496 293 498 295
rect 500 293 508 295
rect 496 289 508 293
rect 520 297 525 306
rect 543 309 557 310
rect 543 307 551 309
rect 553 307 554 309
rect 556 307 557 309
rect 543 306 557 307
rect 567 324 568 326
rect 570 324 572 326
rect 567 319 572 324
rect 567 317 568 319
rect 570 317 572 319
rect 567 315 572 317
rect 543 297 548 306
rect 568 300 572 315
rect 568 298 569 300
rect 571 298 572 300
rect 568 295 572 298
rect 560 293 568 295
rect 570 293 572 295
rect 560 289 572 293
rect 576 326 581 328
rect 576 324 578 326
rect 580 324 581 326
rect 617 333 629 335
rect 617 331 625 333
rect 627 331 629 333
rect 617 329 629 331
rect 576 319 581 324
rect 576 317 578 319
rect 580 317 581 319
rect 576 315 581 317
rect 576 295 580 315
rect 608 320 612 327
rect 617 320 622 329
rect 608 318 622 320
rect 599 317 622 318
rect 599 315 605 317
rect 607 315 619 317
rect 621 315 622 317
rect 599 314 612 315
rect 616 314 622 315
rect 617 313 622 314
rect 591 309 605 310
rect 591 307 595 309
rect 597 307 605 309
rect 591 306 605 307
rect 576 293 578 295
rect 580 293 588 295
rect 576 289 588 293
rect 600 300 605 306
rect 600 298 601 300
rect 603 298 605 300
rect 600 297 605 298
rect 633 304 638 311
rect 661 326 677 327
rect 661 324 663 326
rect 665 324 677 326
rect 661 322 677 324
rect 633 303 635 304
rect 625 302 635 303
rect 637 302 638 304
rect 625 300 638 302
rect 625 298 628 300
rect 630 298 638 300
rect 625 297 638 298
rect 673 294 677 322
rect 653 293 677 294
rect 653 291 655 293
rect 657 291 677 293
rect 653 290 677 291
rect 701 326 706 328
rect 701 324 703 326
rect 705 324 706 326
rect 701 319 706 324
rect 701 317 703 319
rect 705 317 706 319
rect 701 315 706 317
rect 733 326 737 327
rect 733 324 734 326
rect 736 324 737 326
rect 701 295 705 315
rect 733 318 737 324
rect 724 317 737 318
rect 724 315 730 317
rect 732 315 737 317
rect 724 314 737 315
rect 741 318 745 327
rect 772 326 777 328
rect 741 317 754 318
rect 741 315 742 317
rect 744 315 746 317
rect 748 315 754 317
rect 741 314 754 315
rect 716 309 730 310
rect 716 307 717 309
rect 719 307 720 309
rect 722 307 730 309
rect 716 306 730 307
rect 701 293 703 295
rect 705 293 713 295
rect 171 288 195 289
rect 701 289 713 293
rect 725 297 730 306
rect 748 309 762 310
rect 748 307 756 309
rect 758 307 759 309
rect 761 307 762 309
rect 748 306 762 307
rect 772 324 773 326
rect 775 324 777 326
rect 772 319 777 324
rect 772 317 773 319
rect 775 317 777 319
rect 772 315 777 317
rect 748 297 753 306
rect 773 300 777 315
rect 773 298 774 300
rect 776 298 777 300
rect 773 295 777 298
rect 765 293 773 295
rect 775 293 777 295
rect 765 289 777 293
rect 781 326 786 328
rect 781 324 783 326
rect 785 324 786 326
rect 822 333 834 335
rect 822 331 830 333
rect 832 331 834 333
rect 822 329 834 331
rect 781 319 786 324
rect 781 317 783 319
rect 785 317 786 319
rect 781 315 786 317
rect 781 295 785 315
rect 813 320 817 327
rect 822 320 827 329
rect 813 318 827 320
rect 804 317 827 318
rect 804 315 810 317
rect 812 315 824 317
rect 826 315 827 317
rect 804 314 817 315
rect 821 314 827 315
rect 822 313 827 314
rect 796 309 810 310
rect 796 307 800 309
rect 802 307 810 309
rect 796 306 810 307
rect 781 293 783 295
rect 785 293 793 295
rect 781 289 793 293
rect 805 300 810 306
rect 805 298 806 300
rect 808 298 810 300
rect 805 297 810 298
rect 838 304 843 311
rect 866 326 882 327
rect 866 324 868 326
rect 870 324 882 326
rect 866 322 882 324
rect 838 303 840 304
rect 830 302 840 303
rect 842 302 843 304
rect 830 300 843 302
rect 830 298 833 300
rect 835 298 843 300
rect 830 297 843 298
rect 878 294 882 322
rect 1012 297 1210 302
rect 1012 295 1043 297
rect 1045 295 1053 297
rect 1055 295 1083 297
rect 1085 295 1093 297
rect 1095 295 1111 297
rect 1113 295 1164 297
rect 1166 295 1195 297
rect 1197 295 1205 297
rect 1207 295 1210 297
rect 1012 294 1210 295
rect 858 293 882 294
rect 858 291 860 293
rect 862 291 882 293
rect 858 290 882 291
rect 486 283 886 284
rect 4 281 199 282
rect 4 279 17 281
rect 19 279 27 281
rect 29 279 75 281
rect 77 279 85 281
rect 87 279 97 281
rect 99 279 107 281
rect 109 279 138 281
rect 140 279 191 281
rect 193 279 199 281
rect 4 274 199 279
rect 486 281 499 283
rect 501 281 509 283
rect 511 281 557 283
rect 559 281 567 283
rect 569 281 579 283
rect 581 281 589 283
rect 591 281 620 283
rect 622 281 673 283
rect 675 281 704 283
rect 706 281 714 283
rect 716 281 762 283
rect 764 281 772 283
rect 774 281 784 283
rect 786 281 794 283
rect 796 281 825 283
rect 827 281 878 283
rect 880 281 886 283
rect 486 276 886 281
rect 1029 272 1034 281
rect 1046 285 1058 289
rect 1046 283 1054 285
rect 1056 283 1058 285
rect 1054 280 1058 283
rect 1029 271 1043 272
rect 1029 269 1037 271
rect 1039 269 1040 271
rect 1042 269 1043 271
rect 1029 268 1043 269
rect 1022 263 1035 264
rect 1022 261 1027 263
rect 1029 261 1035 263
rect 1022 260 1035 261
rect 1022 255 1026 260
rect 1054 278 1055 280
rect 1057 278 1058 280
rect 1054 263 1058 278
rect 1069 272 1074 281
rect 1086 285 1098 289
rect 1086 283 1094 285
rect 1096 283 1098 285
rect 1069 271 1083 272
rect 1069 269 1077 271
rect 1079 269 1080 271
rect 1082 269 1083 271
rect 1069 268 1083 269
rect 1022 253 1023 255
rect 1025 253 1026 255
rect 1022 251 1026 253
rect 1053 261 1058 263
rect 1053 259 1054 261
rect 1056 259 1058 261
rect 1053 254 1058 259
rect 1053 252 1054 254
rect 1056 252 1058 254
rect 1053 250 1058 252
rect 1062 263 1075 264
rect 1062 261 1067 263
rect 1069 261 1075 263
rect 1062 260 1075 261
rect 1062 256 1066 260
rect 1094 263 1098 283
rect 1062 254 1063 256
rect 1065 254 1066 256
rect 1062 251 1066 254
rect 1093 261 1098 263
rect 1093 259 1094 261
rect 1096 259 1098 261
rect 1093 257 1098 259
rect 1093 255 1094 257
rect 1096 255 1098 257
rect 1093 254 1098 255
rect 1093 252 1094 254
rect 1096 252 1098 254
rect 1093 250 1098 252
rect 1109 287 1133 288
rect 1109 285 1129 287
rect 1131 285 1133 287
rect 1109 284 1133 285
rect 1109 256 1113 284
rect 1148 280 1161 281
rect 1148 278 1156 280
rect 1158 278 1161 280
rect 1148 276 1161 278
rect 1148 274 1149 276
rect 1151 275 1161 276
rect 1151 274 1153 275
rect 1109 254 1125 256
rect 1109 252 1121 254
rect 1123 252 1125 254
rect 1109 251 1125 252
rect 1148 267 1153 274
rect 1181 280 1186 281
rect 1181 278 1183 280
rect 1185 278 1186 280
rect 1181 272 1186 278
rect 1198 285 1210 289
rect 1198 283 1206 285
rect 1208 283 1210 285
rect 1181 271 1195 272
rect 1181 269 1189 271
rect 1191 269 1195 271
rect 1181 268 1195 269
rect 1164 264 1169 265
rect 1164 263 1170 264
rect 1174 263 1187 264
rect 1164 261 1165 263
rect 1167 261 1179 263
rect 1181 261 1187 263
rect 1164 260 1187 261
rect 1164 258 1178 260
rect 1164 249 1169 258
rect 1174 257 1178 258
rect 1206 268 1210 283
rect 1206 266 1207 268
rect 1209 266 1210 268
rect 1206 263 1210 266
rect 1174 255 1175 257
rect 1177 255 1178 257
rect 1174 251 1178 255
rect 1205 261 1210 263
rect 1205 259 1206 261
rect 1208 259 1210 261
rect 1205 254 1210 259
rect 1157 243 1169 249
rect 1205 252 1206 254
rect 1208 252 1210 254
rect 1205 250 1210 252
rect 1021 237 1210 238
rect 1021 235 1053 237
rect 1055 235 1093 237
rect 1095 235 1131 237
rect 1133 235 1205 237
rect 1207 235 1210 237
rect -3 225 1001 230
rect -3 223 4 225
rect 6 223 44 225
rect 46 223 118 225
rect 120 223 149 225
rect 151 223 223 225
rect 225 223 254 225
rect 256 223 294 225
rect 296 223 368 225
rect 370 223 399 225
rect 401 223 473 225
rect 475 223 504 225
rect 506 223 544 225
rect 546 223 618 225
rect 620 223 649 225
rect 651 223 723 225
rect 725 223 754 225
rect 756 223 794 225
rect 796 223 868 225
rect 870 223 899 225
rect 901 223 973 225
rect 975 223 1001 225
rect -3 222 1001 223
rect 1021 225 1210 235
rect 1021 223 1025 225
rect 1027 223 1093 225
rect 1095 223 1105 225
rect 1107 223 1179 225
rect 1181 223 1210 225
rect 1021 222 1210 223
rect 1 216 5 217
rect 1 212 14 216
rect 1 210 3 212
rect 1 205 5 210
rect 1 203 3 205
rect 1 184 5 203
rect 33 208 37 209
rect 33 206 34 208
rect 36 206 37 208
rect 33 200 37 206
rect 16 198 37 200
rect 16 196 30 198
rect 32 196 37 198
rect 41 208 46 210
rect 41 206 43 208
rect 45 206 46 208
rect 82 211 94 217
rect 41 201 46 206
rect 41 199 43 201
rect 45 199 46 201
rect 41 197 46 199
rect 41 192 45 197
rect 1 182 6 184
rect 1 180 3 182
rect 5 180 6 182
rect 1 178 6 180
rect 16 191 45 192
rect 16 189 20 191
rect 22 189 45 191
rect 16 188 45 189
rect 33 179 37 188
rect 41 177 45 188
rect 73 202 77 209
rect 82 202 87 211
rect 73 200 87 202
rect 64 199 87 200
rect 64 197 70 199
rect 72 197 84 199
rect 86 197 87 199
rect 64 196 77 197
rect 81 196 87 197
rect 82 195 87 196
rect 56 191 70 192
rect 56 189 60 191
rect 62 189 70 191
rect 56 188 70 189
rect 41 175 43 177
rect 45 175 53 177
rect 41 171 53 175
rect 65 182 70 188
rect 65 180 66 182
rect 68 180 70 182
rect 65 179 70 180
rect 98 186 103 193
rect 126 208 142 209
rect 126 206 128 208
rect 130 206 142 208
rect 126 204 142 206
rect 98 185 100 186
rect 90 184 100 185
rect 102 184 103 186
rect 90 182 103 184
rect 90 180 93 182
rect 95 180 103 182
rect 90 179 103 180
rect 138 182 142 204
rect 138 180 139 182
rect 141 180 142 182
rect 138 176 142 180
rect 118 175 142 176
rect 118 173 120 175
rect 122 173 142 175
rect 118 172 142 173
rect 146 208 151 210
rect 146 206 148 208
rect 150 206 151 208
rect 187 211 199 217
rect 251 216 255 217
rect 146 201 151 206
rect 146 199 148 201
rect 150 199 151 201
rect 146 197 151 199
rect 146 177 150 197
rect 178 202 182 209
rect 187 202 192 211
rect 251 212 264 216
rect 251 210 253 212
rect 178 200 192 202
rect 169 199 181 200
rect 169 197 175 199
rect 177 198 181 199
rect 183 199 192 200
rect 183 198 189 199
rect 177 197 189 198
rect 191 197 192 199
rect 169 196 182 197
rect 186 196 192 197
rect 187 195 192 196
rect 161 191 175 192
rect 161 189 165 191
rect 167 189 175 191
rect 161 188 175 189
rect 146 175 148 177
rect 150 175 158 177
rect 146 171 158 175
rect 170 182 175 188
rect 170 180 171 182
rect 173 180 175 182
rect 170 179 175 180
rect 203 186 208 193
rect 231 208 247 209
rect 231 206 233 208
rect 235 206 247 208
rect 231 204 247 206
rect 203 185 205 186
rect 195 184 205 185
rect 207 184 208 186
rect 195 182 208 184
rect 195 180 198 182
rect 200 180 208 182
rect 195 179 208 180
rect 243 176 247 204
rect 251 205 255 210
rect 251 203 253 205
rect 251 200 255 203
rect 283 208 287 209
rect 283 206 284 208
rect 286 206 287 208
rect 251 198 252 200
rect 254 198 255 200
rect 251 184 255 198
rect 283 200 287 206
rect 266 198 287 200
rect 266 196 280 198
rect 282 196 287 198
rect 291 208 296 210
rect 291 206 293 208
rect 295 206 296 208
rect 332 211 344 217
rect 291 201 296 206
rect 291 199 293 201
rect 295 199 296 201
rect 291 197 296 199
rect 291 192 295 197
rect 251 182 256 184
rect 251 180 253 182
rect 255 180 256 182
rect 251 178 256 180
rect 266 191 295 192
rect 266 189 270 191
rect 272 189 295 191
rect 266 188 295 189
rect 283 179 287 188
rect 223 175 247 176
rect 223 173 225 175
rect 227 173 247 175
rect 223 172 247 173
rect 291 177 295 188
rect 323 202 327 209
rect 332 202 337 211
rect 323 200 337 202
rect 314 199 337 200
rect 314 197 320 199
rect 322 197 334 199
rect 336 197 337 199
rect 314 196 327 197
rect 331 196 337 197
rect 332 195 337 196
rect 306 191 320 192
rect 306 189 310 191
rect 312 189 320 191
rect 306 188 320 189
rect 291 175 293 177
rect 295 175 303 177
rect 291 171 303 175
rect 315 182 320 188
rect 315 180 316 182
rect 318 180 320 182
rect 315 179 320 180
rect 348 186 353 193
rect 376 208 392 209
rect 376 206 378 208
rect 380 206 392 208
rect 376 204 392 206
rect 348 185 350 186
rect 340 184 350 185
rect 352 184 353 186
rect 340 182 353 184
rect 340 180 343 182
rect 345 180 353 182
rect 340 179 353 180
rect 388 182 392 204
rect 388 180 389 182
rect 391 180 392 182
rect 388 176 392 180
rect 368 175 392 176
rect 368 173 370 175
rect 372 173 392 175
rect 368 172 392 173
rect 396 208 401 210
rect 396 206 398 208
rect 400 206 401 208
rect 437 211 449 217
rect 501 216 505 217
rect 396 201 401 206
rect 396 199 398 201
rect 400 199 401 201
rect 396 197 401 199
rect 396 177 400 197
rect 428 202 432 209
rect 437 202 442 211
rect 501 212 514 216
rect 501 210 503 212
rect 428 200 442 202
rect 419 199 433 200
rect 419 197 425 199
rect 427 198 433 199
rect 435 199 442 200
rect 435 198 439 199
rect 427 197 439 198
rect 441 197 442 199
rect 419 196 432 197
rect 436 196 442 197
rect 437 195 442 196
rect 411 191 425 192
rect 411 189 415 191
rect 417 189 425 191
rect 411 188 425 189
rect 396 175 398 177
rect 400 175 408 177
rect 396 171 408 175
rect 420 182 425 188
rect 420 180 421 182
rect 423 180 425 182
rect 420 179 425 180
rect 453 186 458 193
rect 481 208 497 209
rect 481 206 483 208
rect 485 206 497 208
rect 481 204 497 206
rect 453 185 455 186
rect 445 184 455 185
rect 457 184 458 186
rect 445 182 458 184
rect 445 180 448 182
rect 450 180 458 182
rect 445 179 458 180
rect 493 176 497 204
rect 501 205 505 210
rect 501 203 503 205
rect 501 200 505 203
rect 533 208 537 209
rect 533 206 534 208
rect 536 206 537 208
rect 501 198 502 200
rect 504 198 505 200
rect 501 184 505 198
rect 533 200 537 206
rect 516 198 537 200
rect 516 196 530 198
rect 532 196 537 198
rect 541 208 546 210
rect 541 206 543 208
rect 545 206 546 208
rect 582 211 594 217
rect 541 201 546 206
rect 541 199 543 201
rect 545 199 546 201
rect 541 197 546 199
rect 541 192 545 197
rect 501 182 506 184
rect 501 180 503 182
rect 505 180 506 182
rect 501 178 506 180
rect 516 191 545 192
rect 516 189 520 191
rect 522 189 545 191
rect 516 188 545 189
rect 533 179 537 188
rect 473 175 497 176
rect 473 173 475 175
rect 477 173 497 175
rect 473 172 497 173
rect 541 177 545 188
rect 573 202 577 209
rect 582 202 587 211
rect 573 200 587 202
rect 564 199 587 200
rect 564 197 570 199
rect 572 197 584 199
rect 586 197 587 199
rect 564 196 577 197
rect 581 196 587 197
rect 582 195 587 196
rect 556 191 570 192
rect 556 189 560 191
rect 562 189 570 191
rect 556 188 570 189
rect 541 175 543 177
rect 545 175 553 177
rect 541 171 553 175
rect 565 182 570 188
rect 565 180 566 182
rect 568 180 570 182
rect 565 179 570 180
rect 598 186 603 193
rect 626 208 642 209
rect 626 206 628 208
rect 630 206 642 208
rect 626 204 642 206
rect 598 185 600 186
rect 590 184 600 185
rect 602 184 603 186
rect 590 182 603 184
rect 590 180 593 182
rect 595 180 603 182
rect 590 179 603 180
rect 638 182 642 204
rect 638 180 639 182
rect 641 180 642 182
rect 638 176 642 180
rect 618 175 642 176
rect 618 173 620 175
rect 622 173 642 175
rect 618 172 642 173
rect 646 208 651 210
rect 646 206 648 208
rect 650 206 651 208
rect 687 211 699 217
rect 751 216 755 217
rect 646 201 651 206
rect 646 199 648 201
rect 650 199 651 201
rect 646 197 651 199
rect 646 177 650 197
rect 678 202 682 209
rect 687 202 692 211
rect 751 212 764 216
rect 751 210 753 212
rect 678 200 692 202
rect 669 199 683 200
rect 669 197 675 199
rect 677 198 683 199
rect 685 199 692 200
rect 685 198 689 199
rect 677 197 689 198
rect 691 197 692 199
rect 669 196 682 197
rect 686 196 692 197
rect 687 195 692 196
rect 661 191 675 192
rect 661 189 665 191
rect 667 189 675 191
rect 661 188 675 189
rect 646 175 648 177
rect 650 175 658 177
rect 646 171 658 175
rect 670 182 675 188
rect 670 180 671 182
rect 673 180 675 182
rect 670 179 675 180
rect 703 186 708 193
rect 731 208 747 209
rect 731 206 733 208
rect 735 206 747 208
rect 731 204 747 206
rect 703 185 705 186
rect 695 184 705 185
rect 707 184 708 186
rect 695 182 708 184
rect 695 180 698 182
rect 700 180 708 182
rect 695 179 708 180
rect 743 176 747 204
rect 751 205 755 210
rect 751 203 753 205
rect 751 200 755 203
rect 783 208 787 209
rect 783 206 784 208
rect 786 206 787 208
rect 751 198 752 200
rect 754 198 755 200
rect 751 184 755 198
rect 783 200 787 206
rect 766 198 787 200
rect 766 196 780 198
rect 782 196 787 198
rect 791 208 796 210
rect 791 206 793 208
rect 795 206 796 208
rect 832 211 844 217
rect 791 201 796 206
rect 791 199 793 201
rect 795 199 796 201
rect 791 197 796 199
rect 791 192 795 197
rect 751 182 756 184
rect 751 180 753 182
rect 755 180 756 182
rect 751 178 756 180
rect 766 191 795 192
rect 766 189 770 191
rect 772 189 795 191
rect 766 188 795 189
rect 783 179 787 188
rect 723 175 747 176
rect 723 173 725 175
rect 727 173 747 175
rect 723 172 747 173
rect 791 177 795 188
rect 823 202 827 209
rect 832 202 837 211
rect 823 200 837 202
rect 814 199 837 200
rect 814 197 820 199
rect 822 197 834 199
rect 836 197 837 199
rect 814 196 827 197
rect 831 196 837 197
rect 832 195 837 196
rect 806 191 820 192
rect 806 189 810 191
rect 812 189 820 191
rect 806 188 820 189
rect 791 175 793 177
rect 795 175 803 177
rect 791 171 803 175
rect 815 182 820 188
rect 815 180 816 182
rect 818 180 820 182
rect 815 179 820 180
rect 848 186 853 193
rect 876 208 892 209
rect 876 206 878 208
rect 880 206 892 208
rect 876 204 892 206
rect 848 185 850 186
rect 840 184 850 185
rect 852 184 853 186
rect 840 182 853 184
rect 840 180 843 182
rect 845 180 853 182
rect 840 179 853 180
rect 888 182 892 204
rect 888 180 889 182
rect 891 180 892 182
rect 888 176 892 180
rect 868 175 892 176
rect 868 173 870 175
rect 872 173 892 175
rect 868 172 892 173
rect 896 208 901 210
rect 896 206 898 208
rect 900 206 901 208
rect 937 211 949 217
rect 896 201 901 206
rect 896 199 898 201
rect 900 199 901 201
rect 896 197 901 199
rect 896 177 900 197
rect 928 202 932 209
rect 937 202 942 211
rect 928 200 942 202
rect 919 199 942 200
rect 919 197 925 199
rect 927 197 939 199
rect 941 197 942 199
rect 919 196 932 197
rect 936 196 942 197
rect 937 195 942 196
rect 911 191 925 192
rect 911 189 915 191
rect 917 189 925 191
rect 911 188 925 189
rect 896 175 898 177
rect 900 175 908 177
rect 896 171 908 175
rect 920 182 925 188
rect 920 180 921 182
rect 923 180 925 182
rect 920 179 925 180
rect 953 186 958 193
rect 981 208 997 209
rect 981 206 983 208
rect 985 206 997 208
rect 981 204 997 206
rect 953 185 955 186
rect 945 184 955 185
rect 957 184 958 186
rect 945 182 958 184
rect 945 180 948 182
rect 950 180 958 182
rect 945 179 958 180
rect 993 176 997 204
rect 973 175 997 176
rect 973 173 975 175
rect 977 173 997 175
rect 973 172 997 173
rect 1022 208 1027 210
rect 1022 206 1024 208
rect 1026 206 1027 208
rect 1022 201 1027 206
rect 1022 199 1024 201
rect 1026 199 1027 201
rect 1022 197 1027 199
rect 1054 208 1058 209
rect 1054 206 1055 208
rect 1057 206 1058 208
rect 1022 177 1026 197
rect 1054 200 1058 206
rect 1045 199 1058 200
rect 1045 197 1051 199
rect 1053 197 1058 199
rect 1045 196 1058 197
rect 1062 200 1066 209
rect 1093 208 1098 210
rect 1062 199 1075 200
rect 1062 197 1063 199
rect 1065 197 1067 199
rect 1069 197 1075 199
rect 1062 196 1075 197
rect 1037 191 1051 192
rect 1037 189 1038 191
rect 1040 189 1041 191
rect 1043 189 1051 191
rect 1037 188 1051 189
rect 1022 175 1024 177
rect 1026 175 1034 177
rect 1022 171 1034 175
rect 1046 179 1051 188
rect 1069 191 1083 192
rect 1069 189 1077 191
rect 1079 189 1080 191
rect 1082 189 1083 191
rect 1069 188 1083 189
rect 1093 206 1094 208
rect 1096 206 1098 208
rect 1093 201 1098 206
rect 1093 199 1094 201
rect 1096 199 1098 201
rect 1093 197 1098 199
rect 1069 179 1074 188
rect 1094 182 1098 197
rect 1094 180 1095 182
rect 1097 180 1098 182
rect 1094 177 1098 180
rect 1086 175 1094 177
rect 1096 175 1098 177
rect 1086 171 1098 175
rect 1102 208 1107 210
rect 1102 206 1104 208
rect 1106 206 1107 208
rect 1143 215 1155 217
rect 1143 213 1151 215
rect 1153 213 1155 215
rect 1143 211 1155 213
rect 1102 201 1107 206
rect 1102 199 1104 201
rect 1106 199 1107 201
rect 1102 197 1107 199
rect 1102 177 1106 197
rect 1134 202 1138 209
rect 1143 202 1148 211
rect 1134 200 1148 202
rect 1125 199 1148 200
rect 1125 197 1131 199
rect 1133 197 1145 199
rect 1147 197 1148 199
rect 1125 196 1138 197
rect 1142 196 1148 197
rect 1143 195 1148 196
rect 1117 191 1131 192
rect 1117 189 1121 191
rect 1123 189 1131 191
rect 1117 188 1131 189
rect 1102 175 1104 177
rect 1106 175 1114 177
rect 1102 171 1114 175
rect 1126 182 1131 188
rect 1126 180 1127 182
rect 1129 180 1131 182
rect 1126 179 1131 180
rect 1159 186 1164 193
rect 1187 208 1203 209
rect 1187 206 1189 208
rect 1191 206 1203 208
rect 1187 204 1203 206
rect 1159 185 1161 186
rect 1151 184 1161 185
rect 1163 184 1164 186
rect 1151 182 1164 184
rect 1151 180 1154 182
rect 1156 180 1164 182
rect 1151 179 1164 180
rect 1199 178 1203 204
rect 1199 176 1200 178
rect 1202 176 1203 178
rect 1179 175 1203 176
rect 1179 173 1181 175
rect 1183 173 1203 175
rect 1179 172 1203 173
rect -3 165 1001 166
rect -3 163 4 165
rect 6 163 44 165
rect 46 163 54 165
rect 56 163 85 165
rect 87 163 138 165
rect 140 163 149 165
rect 151 163 159 165
rect 161 163 190 165
rect 192 163 243 165
rect 245 163 254 165
rect 256 163 294 165
rect 296 163 304 165
rect 306 163 335 165
rect 337 163 388 165
rect 390 163 399 165
rect 401 163 409 165
rect 411 163 440 165
rect 442 163 493 165
rect 495 163 504 165
rect 506 163 544 165
rect 546 163 554 165
rect 556 163 585 165
rect 587 163 638 165
rect 640 163 649 165
rect 651 163 659 165
rect 661 163 690 165
rect 692 163 743 165
rect 745 163 754 165
rect 756 163 794 165
rect 796 163 804 165
rect 806 163 835 165
rect 837 163 888 165
rect 890 163 899 165
rect 901 163 909 165
rect 911 163 940 165
rect 942 163 993 165
rect 995 163 1001 165
rect -3 158 1001 163
rect 1012 165 1207 166
rect 1012 163 1025 165
rect 1027 163 1035 165
rect 1037 163 1083 165
rect 1085 163 1093 165
rect 1095 163 1105 165
rect 1107 163 1115 165
rect 1117 163 1146 165
rect 1148 163 1199 165
rect 1201 163 1207 165
rect 1012 158 1207 163
rect 96 145 1215 149
rect 96 144 308 145
rect 96 142 103 144
rect 105 142 113 144
rect 115 142 144 144
rect 146 142 197 144
rect 199 142 218 144
rect 220 142 258 144
rect 260 142 268 144
rect 270 142 299 144
rect 301 143 308 144
rect 310 144 1147 145
rect 310 143 352 144
rect 301 142 352 143
rect 354 142 363 144
rect 365 142 373 144
rect 375 142 404 144
rect 406 142 457 144
rect 459 142 468 144
rect 470 142 508 144
rect 510 142 518 144
rect 520 142 549 144
rect 551 142 558 144
rect 560 142 602 144
rect 604 142 613 144
rect 615 142 623 144
rect 625 142 654 144
rect 656 142 707 144
rect 709 142 718 144
rect 720 142 758 144
rect 760 142 768 144
rect 770 142 799 144
rect 801 142 852 144
rect 854 142 863 144
rect 865 142 873 144
rect 875 142 904 144
rect 906 142 957 144
rect 959 142 968 144
rect 970 142 1008 144
rect 1010 142 1018 144
rect 1020 142 1049 144
rect 1051 142 1102 144
rect 1104 142 1113 144
rect 1115 142 1123 144
rect 1125 143 1147 144
rect 1149 144 1215 145
rect 1149 143 1154 144
rect 1125 142 1154 143
rect 1156 142 1207 144
rect 1209 142 1215 144
rect 96 141 1215 142
rect 100 132 112 136
rect 100 130 102 132
rect 104 130 112 132
rect 177 134 201 135
rect 100 110 104 130
rect 177 132 179 134
rect 181 132 201 134
rect 177 131 201 132
rect 124 127 129 128
rect 124 125 125 127
rect 127 125 129 127
rect 124 119 129 125
rect 100 108 105 110
rect 100 106 102 108
rect 104 106 105 108
rect 100 101 105 106
rect 100 99 102 101
rect 104 99 105 101
rect 115 118 129 119
rect 115 116 116 118
rect 118 116 119 118
rect 121 116 129 118
rect 115 115 129 116
rect 149 127 162 128
rect 149 125 152 127
rect 154 125 162 127
rect 149 123 162 125
rect 149 122 159 123
rect 157 121 159 122
rect 161 121 162 123
rect 141 111 146 112
rect 123 110 146 111
rect 123 108 129 110
rect 131 108 143 110
rect 145 108 146 110
rect 123 107 146 108
rect 132 105 146 107
rect 157 114 162 121
rect 197 113 201 131
rect 255 132 267 136
rect 255 130 257 132
rect 259 130 267 132
rect 332 134 356 135
rect 100 97 105 99
rect 132 98 136 105
rect 141 96 146 105
rect 141 90 153 96
rect 197 111 198 113
rect 200 111 201 113
rect 197 103 201 111
rect 185 101 201 103
rect 185 99 187 101
rect 189 99 201 101
rect 185 98 201 99
rect 215 127 220 129
rect 215 125 217 127
rect 219 125 220 127
rect 215 123 220 125
rect 215 104 219 123
rect 247 119 251 128
rect 255 119 259 130
rect 332 132 334 134
rect 336 132 356 134
rect 332 131 356 132
rect 215 102 217 104
rect 215 97 219 102
rect 215 95 217 97
rect 230 118 259 119
rect 230 116 234 118
rect 236 116 259 118
rect 230 115 259 116
rect 230 109 244 111
rect 246 109 251 111
rect 230 107 251 109
rect 247 101 251 107
rect 247 99 248 101
rect 250 99 251 101
rect 247 98 251 99
rect 255 110 259 115
rect 279 127 284 128
rect 279 125 280 127
rect 282 125 284 127
rect 279 119 284 125
rect 255 108 260 110
rect 255 106 257 108
rect 259 106 260 108
rect 255 101 260 106
rect 255 99 257 101
rect 259 99 260 101
rect 270 118 284 119
rect 270 116 274 118
rect 276 116 284 118
rect 270 115 284 116
rect 304 127 317 128
rect 304 125 307 127
rect 309 125 317 127
rect 304 123 317 125
rect 352 127 356 131
rect 304 122 314 123
rect 312 121 314 122
rect 316 121 317 123
rect 296 111 301 112
rect 278 110 291 111
rect 295 110 301 111
rect 278 108 284 110
rect 286 108 298 110
rect 300 108 301 110
rect 278 107 301 108
rect 287 105 301 107
rect 312 114 317 121
rect 352 125 353 127
rect 355 125 356 127
rect 255 97 260 99
rect 215 91 228 95
rect 215 90 219 91
rect 287 98 291 105
rect 296 96 301 105
rect 296 90 308 96
rect 352 103 356 125
rect 340 101 356 103
rect 340 99 342 101
rect 344 99 356 101
rect 340 98 356 99
rect 360 132 372 136
rect 360 130 362 132
rect 364 130 372 132
rect 437 134 461 135
rect 360 110 364 130
rect 437 132 439 134
rect 441 132 461 134
rect 437 131 461 132
rect 384 127 389 128
rect 384 125 385 127
rect 387 125 389 127
rect 384 119 389 125
rect 360 108 365 110
rect 360 106 362 108
rect 364 106 365 108
rect 360 101 365 106
rect 360 99 362 101
rect 364 99 365 101
rect 375 118 389 119
rect 375 116 379 118
rect 381 116 389 118
rect 375 115 389 116
rect 409 127 422 128
rect 409 125 412 127
rect 414 125 422 127
rect 409 123 422 125
rect 409 122 419 123
rect 417 121 419 122
rect 421 121 422 123
rect 401 111 406 112
rect 383 110 396 111
rect 400 110 406 111
rect 383 108 389 110
rect 391 109 403 110
rect 391 108 395 109
rect 383 107 395 108
rect 397 108 403 109
rect 405 108 406 110
rect 397 107 406 108
rect 392 105 406 107
rect 417 114 422 121
rect 360 97 365 99
rect 392 98 396 105
rect 401 96 406 105
rect 401 90 413 96
rect 457 103 461 131
rect 505 132 517 136
rect 505 130 507 132
rect 509 130 517 132
rect 582 134 606 135
rect 445 101 461 103
rect 445 99 447 101
rect 449 99 458 101
rect 460 99 461 101
rect 445 98 461 99
rect 465 127 470 129
rect 465 125 467 127
rect 469 125 470 127
rect 465 123 470 125
rect 465 109 469 123
rect 465 107 466 109
rect 468 107 469 109
rect 465 104 469 107
rect 497 119 501 128
rect 505 119 509 130
rect 582 132 584 134
rect 586 132 606 134
rect 582 131 606 132
rect 465 102 467 104
rect 465 97 469 102
rect 465 95 467 97
rect 480 118 509 119
rect 480 116 484 118
rect 486 116 509 118
rect 480 115 509 116
rect 480 109 494 111
rect 496 109 501 111
rect 480 107 501 109
rect 497 101 501 107
rect 497 99 498 101
rect 500 99 501 101
rect 497 98 501 99
rect 505 110 509 115
rect 529 127 534 128
rect 529 125 530 127
rect 532 125 534 127
rect 529 119 534 125
rect 505 108 510 110
rect 505 106 507 108
rect 509 106 510 108
rect 505 101 510 106
rect 505 99 507 101
rect 509 99 510 101
rect 520 118 534 119
rect 520 116 524 118
rect 526 116 534 118
rect 520 115 534 116
rect 554 127 567 128
rect 554 125 557 127
rect 559 125 567 127
rect 554 123 567 125
rect 602 127 606 131
rect 554 122 564 123
rect 562 121 564 122
rect 566 121 567 123
rect 546 111 551 112
rect 528 110 541 111
rect 545 110 551 111
rect 528 108 534 110
rect 536 108 548 110
rect 550 108 551 110
rect 528 107 551 108
rect 537 105 551 107
rect 562 114 567 121
rect 602 125 603 127
rect 605 125 606 127
rect 505 97 510 99
rect 465 91 478 95
rect 465 90 469 91
rect 537 98 541 105
rect 546 96 551 105
rect 546 90 558 96
rect 602 103 606 125
rect 590 101 606 103
rect 590 99 592 101
rect 594 99 606 101
rect 590 98 606 99
rect 610 132 622 136
rect 610 130 612 132
rect 614 130 622 132
rect 687 134 711 135
rect 610 110 614 130
rect 687 132 689 134
rect 691 132 711 134
rect 687 131 711 132
rect 634 127 639 128
rect 634 125 635 127
rect 637 125 639 127
rect 634 119 639 125
rect 610 108 615 110
rect 610 106 612 108
rect 614 106 615 108
rect 610 101 615 106
rect 610 99 612 101
rect 614 99 615 101
rect 625 118 639 119
rect 625 116 629 118
rect 631 116 639 118
rect 625 115 639 116
rect 659 127 672 128
rect 659 125 662 127
rect 664 125 672 127
rect 659 123 672 125
rect 659 122 669 123
rect 667 121 669 122
rect 671 121 672 123
rect 651 111 656 112
rect 633 110 646 111
rect 650 110 656 111
rect 633 108 639 110
rect 641 109 653 110
rect 641 108 647 109
rect 633 107 647 108
rect 649 108 653 109
rect 655 108 656 110
rect 649 107 656 108
rect 642 105 656 107
rect 667 114 672 121
rect 610 97 615 99
rect 642 98 646 105
rect 651 96 656 105
rect 651 90 663 96
rect 707 103 711 131
rect 755 132 767 136
rect 755 130 757 132
rect 759 130 767 132
rect 832 134 856 135
rect 695 101 711 103
rect 695 99 697 101
rect 699 99 708 101
rect 710 99 711 101
rect 695 98 711 99
rect 715 127 720 129
rect 715 125 717 127
rect 719 125 720 127
rect 715 123 720 125
rect 715 109 719 123
rect 715 107 716 109
rect 718 107 719 109
rect 715 104 719 107
rect 747 119 751 128
rect 755 119 759 130
rect 832 132 834 134
rect 836 132 856 134
rect 832 131 856 132
rect 715 102 717 104
rect 715 97 719 102
rect 715 95 717 97
rect 730 118 759 119
rect 730 116 734 118
rect 736 116 759 118
rect 730 115 759 116
rect 730 109 744 111
rect 746 109 751 111
rect 730 107 751 109
rect 747 101 751 107
rect 747 99 748 101
rect 750 99 751 101
rect 747 98 751 99
rect 755 110 759 115
rect 779 127 784 128
rect 779 125 780 127
rect 782 125 784 127
rect 779 119 784 125
rect 755 108 760 110
rect 755 106 757 108
rect 759 106 760 108
rect 755 101 760 106
rect 755 99 757 101
rect 759 99 760 101
rect 770 118 784 119
rect 770 116 774 118
rect 776 116 784 118
rect 770 115 784 116
rect 804 127 817 128
rect 804 125 807 127
rect 809 125 817 127
rect 804 123 817 125
rect 852 127 856 131
rect 804 122 814 123
rect 812 121 814 122
rect 816 121 817 123
rect 796 111 801 112
rect 778 110 791 111
rect 795 110 801 111
rect 778 108 784 110
rect 786 108 798 110
rect 800 108 801 110
rect 778 107 801 108
rect 787 105 801 107
rect 812 114 817 121
rect 852 125 853 127
rect 855 125 856 127
rect 755 97 760 99
rect 715 91 728 95
rect 715 90 719 91
rect 787 98 791 105
rect 796 96 801 105
rect 796 90 808 96
rect 852 103 856 125
rect 840 101 856 103
rect 840 99 842 101
rect 844 99 856 101
rect 840 98 856 99
rect 860 132 872 136
rect 860 130 862 132
rect 864 130 872 132
rect 937 134 961 135
rect 860 110 864 130
rect 937 132 939 134
rect 941 132 961 134
rect 937 131 961 132
rect 884 127 889 128
rect 884 125 885 127
rect 887 125 889 127
rect 884 119 889 125
rect 860 108 865 110
rect 860 106 862 108
rect 864 106 865 108
rect 860 101 865 106
rect 860 99 862 101
rect 864 99 865 101
rect 875 118 889 119
rect 875 116 879 118
rect 881 116 889 118
rect 875 115 889 116
rect 909 127 922 128
rect 909 125 912 127
rect 914 125 922 127
rect 909 123 922 125
rect 909 122 919 123
rect 917 121 919 122
rect 921 121 922 123
rect 901 111 906 112
rect 883 110 896 111
rect 900 110 906 111
rect 883 108 889 110
rect 891 109 903 110
rect 891 108 897 109
rect 883 107 897 108
rect 899 108 903 109
rect 905 108 906 110
rect 899 107 906 108
rect 892 105 906 107
rect 917 114 922 121
rect 860 97 865 99
rect 892 98 896 105
rect 901 96 906 105
rect 901 90 913 96
rect 957 103 961 131
rect 1005 132 1017 136
rect 1005 130 1007 132
rect 1009 130 1017 132
rect 1082 134 1106 135
rect 945 101 961 103
rect 945 99 947 101
rect 949 99 961 101
rect 945 98 961 99
rect 965 127 970 129
rect 965 125 967 127
rect 969 125 970 127
rect 965 123 970 125
rect 965 109 969 123
rect 965 107 966 109
rect 968 107 969 109
rect 965 104 969 107
rect 997 119 1001 128
rect 1005 119 1009 130
rect 1082 132 1084 134
rect 1086 132 1106 134
rect 1082 131 1106 132
rect 965 102 967 104
rect 965 97 969 102
rect 965 95 967 97
rect 980 118 1009 119
rect 980 116 984 118
rect 986 116 1009 118
rect 980 115 1009 116
rect 980 109 994 111
rect 996 109 1001 111
rect 980 107 1001 109
rect 997 101 1001 107
rect 997 99 998 101
rect 1000 99 1001 101
rect 997 98 1001 99
rect 1005 110 1009 115
rect 1029 127 1034 128
rect 1029 125 1030 127
rect 1032 125 1034 127
rect 1029 119 1034 125
rect 1005 108 1010 110
rect 1005 106 1007 108
rect 1009 106 1010 108
rect 1005 101 1010 106
rect 1005 99 1007 101
rect 1009 99 1010 101
rect 1020 118 1034 119
rect 1020 116 1024 118
rect 1026 116 1034 118
rect 1020 115 1034 116
rect 1054 127 1067 128
rect 1054 125 1057 127
rect 1059 125 1067 127
rect 1054 123 1067 125
rect 1102 127 1106 131
rect 1054 122 1064 123
rect 1062 121 1064 122
rect 1066 121 1067 123
rect 1046 111 1051 112
rect 1028 110 1041 111
rect 1045 110 1051 111
rect 1028 108 1034 110
rect 1036 108 1048 110
rect 1050 108 1051 110
rect 1028 107 1051 108
rect 1037 105 1051 107
rect 1062 114 1067 121
rect 1102 125 1103 127
rect 1105 125 1106 127
rect 1005 97 1010 99
rect 965 91 978 95
rect 965 90 969 91
rect 1037 98 1041 105
rect 1046 96 1051 105
rect 1046 90 1058 96
rect 1102 103 1106 125
rect 1090 101 1106 103
rect 1090 99 1092 101
rect 1094 99 1106 101
rect 1090 98 1106 99
rect 1110 132 1122 136
rect 1110 130 1112 132
rect 1114 130 1122 132
rect 1187 134 1211 135
rect 1110 110 1114 130
rect 1187 132 1189 134
rect 1191 132 1211 134
rect 1187 131 1211 132
rect 1134 127 1139 128
rect 1134 125 1135 127
rect 1137 125 1139 127
rect 1134 119 1139 125
rect 1110 108 1115 110
rect 1110 106 1112 108
rect 1114 106 1115 108
rect 1110 101 1115 106
rect 1110 99 1112 101
rect 1114 99 1115 101
rect 1125 118 1139 119
rect 1125 116 1129 118
rect 1131 116 1139 118
rect 1125 115 1139 116
rect 1159 127 1172 128
rect 1159 125 1162 127
rect 1164 125 1172 127
rect 1159 123 1172 125
rect 1159 122 1169 123
rect 1167 121 1169 122
rect 1171 121 1172 123
rect 1151 111 1156 112
rect 1133 110 1156 111
rect 1133 108 1139 110
rect 1141 108 1147 110
rect 1149 108 1153 110
rect 1155 108 1156 110
rect 1133 107 1156 108
rect 1142 105 1156 107
rect 1167 114 1172 121
rect 1110 97 1115 99
rect 1142 98 1146 105
rect 1151 96 1156 105
rect 1151 90 1163 96
rect 1207 103 1211 131
rect 1195 101 1211 103
rect 1195 99 1197 101
rect 1199 99 1211 101
rect 1195 98 1211 99
rect 96 84 1215 85
rect 96 82 103 84
rect 105 82 177 84
rect 179 82 218 84
rect 220 82 258 84
rect 260 82 332 84
rect 334 82 363 84
rect 365 82 437 84
rect 439 82 468 84
rect 470 82 508 84
rect 510 82 582 84
rect 584 82 613 84
rect 615 82 687 84
rect 689 82 718 84
rect 720 82 758 84
rect 760 82 832 84
rect 834 82 863 84
rect 865 82 937 84
rect 939 82 968 84
rect 970 82 1008 84
rect 1010 82 1082 84
rect 1084 82 1113 84
rect 1115 82 1187 84
rect 1189 82 1215 84
rect 96 77 1215 82
rect 3 72 1012 77
rect 3 70 10 72
rect 12 70 50 72
rect 52 70 124 72
rect 126 70 155 72
rect 157 70 229 72
rect 231 70 260 72
rect 262 70 300 72
rect 302 70 374 72
rect 376 70 405 72
rect 407 70 479 72
rect 481 70 510 72
rect 512 70 550 72
rect 552 70 624 72
rect 626 70 655 72
rect 657 70 729 72
rect 731 70 760 72
rect 762 70 800 72
rect 802 70 874 72
rect 876 70 905 72
rect 907 70 979 72
rect 981 71 1012 72
rect 981 70 1007 71
rect 3 69 1007 70
rect 7 63 11 64
rect 7 59 20 63
rect 7 57 9 59
rect 7 52 11 57
rect 7 50 9 52
rect 7 31 11 50
rect 39 55 43 56
rect 39 53 40 55
rect 42 53 43 55
rect 39 47 43 53
rect 22 45 43 47
rect 22 43 36 45
rect 38 43 43 45
rect 47 55 52 57
rect 47 53 49 55
rect 51 53 52 55
rect 88 58 100 64
rect 47 48 52 53
rect 47 46 49 48
rect 51 46 52 48
rect 47 44 52 46
rect 47 39 51 44
rect 7 29 12 31
rect 7 27 9 29
rect 11 27 12 29
rect 7 25 12 27
rect 22 38 51 39
rect 22 36 26 38
rect 28 36 51 38
rect 22 35 51 36
rect 39 26 43 35
rect 47 24 51 35
rect 79 49 83 56
rect 88 49 93 58
rect 79 47 93 49
rect 70 46 93 47
rect 70 44 76 46
rect 78 44 90 46
rect 92 44 93 46
rect 70 43 83 44
rect 87 43 93 44
rect 88 42 93 43
rect 62 38 76 39
rect 62 36 66 38
rect 68 36 76 38
rect 62 35 76 36
rect 47 22 49 24
rect 51 22 59 24
rect 47 18 59 22
rect 71 29 76 35
rect 71 27 72 29
rect 74 27 76 29
rect 71 26 76 27
rect 104 38 109 40
rect 104 36 106 38
rect 108 36 109 38
rect 104 33 109 36
rect 132 55 148 56
rect 132 53 134 55
rect 136 53 148 55
rect 132 51 148 53
rect 104 32 106 33
rect 96 31 106 32
rect 108 31 109 33
rect 96 29 109 31
rect 96 27 99 29
rect 101 27 109 29
rect 96 26 109 27
rect 144 29 148 51
rect 144 27 145 29
rect 147 27 148 29
rect 144 23 148 27
rect 124 22 148 23
rect 124 20 126 22
rect 128 20 148 22
rect 124 19 148 20
rect 152 55 157 57
rect 152 53 154 55
rect 156 53 157 55
rect 193 58 205 64
rect 257 63 261 64
rect 152 48 157 53
rect 152 46 154 48
rect 156 46 157 48
rect 152 44 157 46
rect 152 24 156 44
rect 184 49 188 56
rect 193 49 198 58
rect 257 59 270 63
rect 257 57 259 59
rect 184 47 198 49
rect 175 46 187 47
rect 175 44 181 46
rect 183 45 187 46
rect 189 46 198 47
rect 189 45 195 46
rect 183 44 195 45
rect 197 44 198 46
rect 175 43 188 44
rect 192 43 198 44
rect 193 42 198 43
rect 167 38 181 39
rect 167 36 171 38
rect 173 36 181 38
rect 167 35 181 36
rect 152 22 154 24
rect 156 22 164 24
rect 152 18 164 22
rect 176 29 181 35
rect 176 27 177 29
rect 179 27 181 29
rect 176 26 181 27
rect 209 33 214 40
rect 237 55 253 56
rect 237 53 239 55
rect 241 53 253 55
rect 237 51 253 53
rect 209 32 211 33
rect 201 31 211 32
rect 213 31 214 33
rect 201 29 214 31
rect 201 27 204 29
rect 206 27 214 29
rect 201 26 214 27
rect 249 23 253 51
rect 257 52 261 57
rect 257 50 259 52
rect 257 47 261 50
rect 289 55 293 56
rect 289 53 290 55
rect 292 53 293 55
rect 257 45 258 47
rect 260 45 261 47
rect 257 31 261 45
rect 289 47 293 53
rect 272 45 293 47
rect 272 43 286 45
rect 288 43 293 45
rect 297 55 302 57
rect 297 53 299 55
rect 301 53 302 55
rect 338 58 350 64
rect 297 48 302 53
rect 297 46 299 48
rect 301 46 302 48
rect 297 44 302 46
rect 297 39 301 44
rect 257 29 262 31
rect 257 27 259 29
rect 261 27 262 29
rect 257 25 262 27
rect 272 38 301 39
rect 272 36 276 38
rect 278 36 301 38
rect 272 35 301 36
rect 289 26 293 35
rect 229 22 253 23
rect 229 20 231 22
rect 233 20 253 22
rect 229 19 253 20
rect 297 24 301 35
rect 329 49 333 56
rect 338 49 343 58
rect 329 47 343 49
rect 320 46 343 47
rect 320 44 326 46
rect 328 44 340 46
rect 342 44 343 46
rect 320 43 333 44
rect 337 43 343 44
rect 338 42 343 43
rect 312 38 326 39
rect 312 36 316 38
rect 318 36 326 38
rect 312 35 326 36
rect 297 22 299 24
rect 301 22 309 24
rect 297 18 309 22
rect 321 29 326 35
rect 321 27 322 29
rect 324 27 326 29
rect 321 26 326 27
rect 354 39 359 40
rect 354 37 356 39
rect 358 37 359 39
rect 354 33 359 37
rect 382 55 398 56
rect 382 53 384 55
rect 386 53 398 55
rect 382 51 398 53
rect 354 32 356 33
rect 346 31 356 32
rect 358 31 359 33
rect 346 29 359 31
rect 346 27 349 29
rect 351 27 359 29
rect 346 26 359 27
rect 394 29 398 51
rect 394 27 395 29
rect 397 27 398 29
rect 394 23 398 27
rect 374 22 398 23
rect 374 20 376 22
rect 378 20 398 22
rect 374 19 398 20
rect 402 55 407 57
rect 402 53 404 55
rect 406 53 407 55
rect 443 58 455 64
rect 507 63 511 64
rect 402 48 407 53
rect 402 46 404 48
rect 406 46 407 48
rect 402 44 407 46
rect 402 24 406 44
rect 434 49 438 56
rect 443 49 448 58
rect 507 59 520 63
rect 507 57 509 59
rect 434 47 448 49
rect 425 46 439 47
rect 425 44 431 46
rect 433 45 439 46
rect 441 46 448 47
rect 441 45 445 46
rect 433 44 445 45
rect 447 44 448 46
rect 425 43 438 44
rect 442 43 448 44
rect 443 42 448 43
rect 417 38 431 39
rect 417 36 421 38
rect 423 36 431 38
rect 417 35 431 36
rect 402 22 404 24
rect 406 22 414 24
rect 402 18 414 22
rect 426 29 431 35
rect 426 27 427 29
rect 429 27 431 29
rect 426 26 431 27
rect 459 33 464 40
rect 487 55 503 56
rect 487 53 489 55
rect 491 53 503 55
rect 487 51 503 53
rect 459 32 461 33
rect 451 31 461 32
rect 463 31 464 33
rect 451 29 464 31
rect 451 27 454 29
rect 456 27 464 29
rect 451 26 464 27
rect 499 23 503 51
rect 507 52 511 57
rect 507 50 509 52
rect 507 47 511 50
rect 539 55 543 56
rect 539 53 540 55
rect 542 53 543 55
rect 507 45 508 47
rect 510 45 511 47
rect 507 31 511 45
rect 539 47 543 53
rect 522 45 543 47
rect 522 43 536 45
rect 538 43 543 45
rect 547 55 552 57
rect 547 53 549 55
rect 551 53 552 55
rect 588 58 600 64
rect 547 48 552 53
rect 547 46 549 48
rect 551 46 552 48
rect 547 44 552 46
rect 547 39 551 44
rect 507 29 512 31
rect 507 27 509 29
rect 511 27 512 29
rect 507 25 512 27
rect 522 38 551 39
rect 522 36 526 38
rect 528 36 551 38
rect 522 35 551 36
rect 539 26 543 35
rect 479 22 503 23
rect 479 20 481 22
rect 483 20 503 22
rect 479 19 503 20
rect 547 24 551 35
rect 579 49 583 56
rect 588 49 593 58
rect 579 47 593 49
rect 570 46 593 47
rect 570 44 576 46
rect 578 44 590 46
rect 592 44 593 46
rect 570 43 583 44
rect 587 43 593 44
rect 588 42 593 43
rect 562 38 576 39
rect 562 36 566 38
rect 568 36 576 38
rect 562 35 576 36
rect 547 22 549 24
rect 551 22 559 24
rect 547 18 559 22
rect 571 29 576 35
rect 571 27 572 29
rect 574 27 576 29
rect 571 26 576 27
rect 604 39 609 40
rect 604 37 606 39
rect 608 37 609 39
rect 604 33 609 37
rect 632 55 648 56
rect 632 53 634 55
rect 636 53 648 55
rect 632 51 648 53
rect 604 32 606 33
rect 596 31 606 32
rect 608 31 609 33
rect 596 29 609 31
rect 596 27 599 29
rect 601 27 609 29
rect 596 26 609 27
rect 644 29 648 51
rect 644 27 645 29
rect 647 27 648 29
rect 644 23 648 27
rect 624 22 648 23
rect 624 20 626 22
rect 628 20 648 22
rect 624 19 648 20
rect 652 55 657 57
rect 652 53 654 55
rect 656 53 657 55
rect 693 58 705 64
rect 757 63 761 64
rect 652 48 657 53
rect 652 46 654 48
rect 656 46 657 48
rect 652 44 657 46
rect 652 24 656 44
rect 684 49 688 56
rect 693 49 698 58
rect 757 59 770 63
rect 757 57 759 59
rect 684 47 698 49
rect 675 46 689 47
rect 675 44 681 46
rect 683 45 689 46
rect 691 46 698 47
rect 691 45 695 46
rect 683 44 695 45
rect 697 44 698 46
rect 675 43 688 44
rect 692 43 698 44
rect 693 42 698 43
rect 667 38 681 39
rect 667 36 671 38
rect 673 36 681 38
rect 667 35 681 36
rect 652 22 654 24
rect 656 22 664 24
rect 652 18 664 22
rect 676 29 681 35
rect 676 27 677 29
rect 679 27 681 29
rect 676 26 681 27
rect 709 33 714 40
rect 737 55 753 56
rect 737 53 739 55
rect 741 53 753 55
rect 737 51 753 53
rect 709 32 711 33
rect 701 31 711 32
rect 713 31 714 33
rect 701 29 714 31
rect 701 27 704 29
rect 706 27 714 29
rect 701 26 714 27
rect 749 23 753 51
rect 757 52 761 57
rect 757 50 759 52
rect 757 47 761 50
rect 789 55 793 56
rect 789 53 790 55
rect 792 53 793 55
rect 757 45 758 47
rect 760 45 761 47
rect 757 31 761 45
rect 789 47 793 53
rect 772 45 793 47
rect 772 43 786 45
rect 788 43 793 45
rect 797 55 802 57
rect 797 53 799 55
rect 801 53 802 55
rect 838 58 850 64
rect 797 48 802 53
rect 797 46 799 48
rect 801 46 802 48
rect 797 44 802 46
rect 797 39 801 44
rect 757 29 762 31
rect 757 27 759 29
rect 761 27 762 29
rect 757 25 762 27
rect 772 38 801 39
rect 772 36 776 38
rect 778 36 801 38
rect 772 35 801 36
rect 789 26 793 35
rect 729 22 753 23
rect 729 20 731 22
rect 733 20 753 22
rect 729 19 753 20
rect 797 24 801 35
rect 829 49 833 56
rect 838 49 843 58
rect 829 47 843 49
rect 820 46 843 47
rect 820 44 826 46
rect 828 44 840 46
rect 842 44 843 46
rect 820 43 833 44
rect 837 43 843 44
rect 838 42 843 43
rect 812 38 826 39
rect 812 36 816 38
rect 818 36 826 38
rect 812 35 826 36
rect 797 22 799 24
rect 801 22 809 24
rect 797 18 809 22
rect 821 29 826 35
rect 821 27 822 29
rect 824 27 826 29
rect 821 26 826 27
rect 854 38 859 40
rect 854 36 856 38
rect 858 36 859 38
rect 854 33 859 36
rect 882 55 898 56
rect 882 53 884 55
rect 886 53 898 55
rect 882 51 898 53
rect 854 32 856 33
rect 846 31 856 32
rect 858 31 859 33
rect 846 29 859 31
rect 846 27 849 29
rect 851 27 859 29
rect 846 26 859 27
rect 894 29 898 51
rect 894 27 895 29
rect 897 27 898 29
rect 894 23 898 27
rect 874 22 898 23
rect 874 20 876 22
rect 878 20 898 22
rect 874 19 898 20
rect 902 55 907 57
rect 902 53 904 55
rect 906 53 907 55
rect 943 58 955 64
rect 902 48 907 53
rect 902 46 904 48
rect 906 46 907 48
rect 902 44 907 46
rect 902 24 906 44
rect 934 49 938 56
rect 943 49 948 58
rect 934 47 948 49
rect 925 46 948 47
rect 925 44 931 46
rect 933 44 939 46
rect 941 44 945 46
rect 947 44 948 46
rect 925 43 948 44
rect 943 42 948 43
rect 917 38 931 39
rect 917 36 921 38
rect 923 36 931 38
rect 917 35 931 36
rect 902 22 904 24
rect 906 22 914 24
rect 902 18 914 22
rect 926 29 931 35
rect 926 27 927 29
rect 929 27 931 29
rect 926 26 931 27
rect 959 33 964 40
rect 987 55 1003 56
rect 987 53 989 55
rect 991 53 1003 55
rect 987 51 1003 53
rect 959 32 961 33
rect 951 31 961 32
rect 963 31 964 33
rect 951 29 964 31
rect 951 27 954 29
rect 956 27 964 29
rect 951 26 964 27
rect 999 23 1003 51
rect 979 22 1003 23
rect 979 20 981 22
rect 983 20 1003 22
rect 979 19 1003 20
rect 3 12 1007 13
rect 3 10 10 12
rect 12 10 50 12
rect 52 10 60 12
rect 62 10 91 12
rect 93 10 144 12
rect 146 10 155 12
rect 157 10 165 12
rect 167 10 196 12
rect 198 10 249 12
rect 251 10 260 12
rect 262 10 300 12
rect 302 10 310 12
rect 312 10 341 12
rect 343 10 394 12
rect 396 10 405 12
rect 407 10 415 12
rect 417 10 446 12
rect 448 10 499 12
rect 501 10 510 12
rect 512 10 550 12
rect 552 10 560 12
rect 562 10 591 12
rect 593 10 644 12
rect 646 10 655 12
rect 657 10 665 12
rect 667 10 696 12
rect 698 10 749 12
rect 751 10 760 12
rect 762 10 800 12
rect 802 10 810 12
rect 812 10 841 12
rect 843 10 894 12
rect 896 10 905 12
rect 907 10 915 12
rect 917 11 946 12
rect 917 10 939 11
rect 3 9 939 10
rect 941 10 946 11
rect 948 10 999 12
rect 1001 10 1007 12
rect 941 9 1007 10
rect 3 5 1007 9
<< alu2 >>
rect 528 398 660 399
rect 46 396 178 397
rect 46 394 47 396
rect 49 394 148 396
rect 150 394 175 396
rect 177 394 178 396
rect 528 396 529 398
rect 531 396 630 398
rect 632 396 657 398
rect 659 396 660 398
rect 528 395 660 396
rect 733 398 865 399
rect 733 396 734 398
rect 736 396 835 398
rect 837 396 862 398
rect 864 396 865 398
rect 733 395 865 396
rect 46 393 178 394
rect 511 389 517 390
rect 29 387 35 388
rect 29 385 32 387
rect 34 385 35 387
rect 6 371 18 372
rect 6 369 15 371
rect 17 369 18 371
rect 6 367 18 369
rect 6 294 11 367
rect 29 307 35 385
rect 71 387 75 388
rect 71 385 72 387
rect 74 385 75 387
rect 54 372 58 373
rect 54 370 55 372
rect 57 370 58 372
rect 54 346 58 370
rect 46 342 58 346
rect 46 324 50 342
rect 46 322 47 324
rect 49 322 50 324
rect 46 321 50 322
rect 29 305 30 307
rect 32 305 35 307
rect 29 304 35 305
rect 54 315 58 316
rect 54 313 55 315
rect 57 313 58 315
rect 54 294 58 313
rect 71 307 75 385
rect 198 384 202 388
rect 198 382 199 384
rect 201 382 202 384
rect 85 373 170 374
rect 85 371 86 373
rect 88 371 167 373
rect 169 371 170 373
rect 85 370 170 371
rect 198 347 202 382
rect 511 387 514 389
rect 516 387 517 389
rect 142 342 202 347
rect 488 373 500 374
rect 488 371 497 373
rect 499 371 500 373
rect 488 369 500 371
rect 142 331 147 342
rect 142 329 143 331
rect 145 329 147 331
rect 142 327 147 329
rect 71 305 72 307
rect 74 305 75 307
rect 71 304 75 305
rect 86 298 151 299
rect 86 296 87 298
rect 89 296 119 298
rect 121 296 146 298
rect 148 296 151 298
rect 86 295 151 296
rect 488 296 493 369
rect 511 309 517 387
rect 553 389 557 390
rect 553 387 554 389
rect 556 387 557 389
rect 536 374 540 375
rect 536 372 537 374
rect 539 372 540 374
rect 536 348 540 372
rect 528 344 540 348
rect 528 326 532 344
rect 528 324 529 326
rect 531 324 532 326
rect 528 323 532 324
rect 511 307 512 309
rect 514 307 517 309
rect 511 306 517 307
rect 536 317 540 318
rect 536 315 537 317
rect 539 315 540 317
rect 536 296 540 315
rect 553 309 557 387
rect 680 386 684 390
rect 680 384 681 386
rect 683 384 684 386
rect 567 375 652 376
rect 567 373 568 375
rect 570 373 649 375
rect 651 373 652 375
rect 567 372 652 373
rect 680 349 684 384
rect 716 389 722 390
rect 716 387 719 389
rect 721 387 722 389
rect 624 344 684 349
rect 693 373 705 374
rect 693 371 702 373
rect 704 371 705 373
rect 693 369 705 371
rect 624 333 629 344
rect 624 331 625 333
rect 627 331 629 333
rect 624 329 629 331
rect 553 307 554 309
rect 556 307 557 309
rect 553 306 557 307
rect 568 300 633 301
rect 568 298 569 300
rect 571 298 601 300
rect 603 298 628 300
rect 630 298 633 300
rect 568 297 633 298
rect 568 296 606 297
rect 693 296 698 369
rect 716 309 722 387
rect 758 389 762 390
rect 758 387 759 389
rect 761 387 762 389
rect 741 374 745 375
rect 741 372 742 374
rect 744 372 745 374
rect 741 348 745 372
rect 733 344 745 348
rect 733 326 737 344
rect 733 324 734 326
rect 736 324 737 326
rect 733 323 737 324
rect 716 307 717 309
rect 719 307 722 309
rect 716 306 722 307
rect 741 317 745 318
rect 741 315 742 317
rect 744 315 745 317
rect 741 296 745 315
rect 758 309 762 387
rect 885 386 889 390
rect 885 384 886 386
rect 888 384 889 386
rect 772 375 857 376
rect 772 373 773 375
rect 775 373 854 375
rect 856 373 857 375
rect 772 372 857 373
rect 885 349 889 384
rect 829 344 889 349
rect 829 333 834 344
rect 829 331 830 333
rect 832 331 834 333
rect 829 329 834 331
rect 758 307 759 309
rect 761 307 762 309
rect 758 306 762 307
rect 773 300 838 301
rect 773 298 774 300
rect 776 298 806 300
rect 808 298 833 300
rect 835 298 838 300
rect 773 297 838 298
rect 773 296 811 297
rect 86 294 124 295
rect 6 290 58 294
rect 488 292 540 296
rect 693 292 745 296
rect 1054 280 1186 281
rect 1054 278 1055 280
rect 1057 278 1156 280
rect 1158 278 1183 280
rect 1185 278 1186 280
rect 1054 277 1186 278
rect 1037 271 1043 272
rect 1037 269 1040 271
rect 1042 269 1043 271
rect 1014 255 1026 256
rect 1014 253 1023 255
rect 1025 253 1026 255
rect 1014 251 1026 253
rect 33 208 151 209
rect 33 206 34 208
rect 36 206 148 208
rect 150 206 151 208
rect 33 205 151 206
rect 283 208 401 209
rect 283 206 284 208
rect 286 206 398 208
rect 400 206 401 208
rect 283 205 401 206
rect 533 208 651 209
rect 533 206 534 208
rect 536 206 648 208
rect 650 206 651 208
rect 533 205 651 206
rect 783 208 901 209
rect 783 206 784 208
rect 786 206 898 208
rect 900 206 901 208
rect 783 205 901 206
rect 180 200 255 201
rect 180 198 181 200
rect 183 198 252 200
rect 254 198 255 200
rect 180 197 255 198
rect 432 200 505 201
rect 432 198 433 200
rect 435 198 502 200
rect 504 198 505 200
rect 432 197 505 198
rect 682 200 755 201
rect 682 198 683 200
rect 685 198 752 200
rect 754 198 755 200
rect 682 197 755 198
rect 1 182 6 184
rect 1 180 3 182
rect 5 180 6 182
rect 1 178 6 180
rect 65 182 98 183
rect 65 180 66 182
rect 68 180 93 182
rect 95 180 98 182
rect 65 179 98 180
rect 138 182 203 183
rect 138 180 139 182
rect 141 180 171 182
rect 173 180 198 182
rect 200 180 203 182
rect 138 179 203 180
rect 315 182 348 183
rect 315 180 316 182
rect 318 180 343 182
rect 345 180 348 182
rect 315 179 348 180
rect 388 182 453 183
rect 388 180 389 182
rect 391 180 421 182
rect 423 180 448 182
rect 450 180 453 182
rect 388 179 453 180
rect 565 182 598 183
rect 565 180 566 182
rect 568 180 593 182
rect 595 180 598 182
rect 565 179 598 180
rect 638 182 703 183
rect 638 180 639 182
rect 641 180 671 182
rect 673 180 698 182
rect 700 180 703 182
rect 638 179 703 180
rect 815 182 848 183
rect 815 180 816 182
rect 818 180 843 182
rect 845 180 848 182
rect 815 179 848 180
rect 888 182 953 183
rect 888 180 889 182
rect 891 180 921 182
rect 923 180 948 182
rect 950 180 953 182
rect 888 179 953 180
rect 1014 178 1019 251
rect 1037 191 1043 269
rect 1079 271 1083 272
rect 1079 269 1080 271
rect 1082 269 1083 271
rect 1062 256 1066 257
rect 1062 254 1063 256
rect 1065 254 1066 256
rect 1062 230 1066 254
rect 1054 226 1066 230
rect 1054 208 1058 226
rect 1054 206 1055 208
rect 1057 206 1058 208
rect 1054 205 1058 206
rect 1037 189 1038 191
rect 1040 189 1043 191
rect 1037 188 1043 189
rect 1062 199 1066 200
rect 1062 197 1063 199
rect 1065 197 1066 199
rect 1062 178 1066 197
rect 1079 191 1083 269
rect 1206 268 1210 272
rect 1206 266 1207 268
rect 1209 266 1210 268
rect 1093 257 1178 258
rect 1093 255 1094 257
rect 1096 255 1175 257
rect 1177 255 1178 257
rect 1093 254 1178 255
rect 1206 231 1210 266
rect 1150 226 1210 231
rect 1150 215 1155 226
rect 1150 213 1151 215
rect 1153 213 1155 215
rect 1150 211 1155 213
rect 1079 189 1080 191
rect 1082 189 1083 191
rect 1079 188 1083 189
rect 1102 190 1106 191
rect 1102 188 1103 190
rect 1105 188 1106 190
rect 1102 187 1106 188
rect 1094 182 1159 183
rect 1094 180 1095 182
rect 1097 180 1127 182
rect 1129 180 1154 182
rect 1156 180 1159 182
rect 1094 179 1159 180
rect 1094 178 1132 179
rect 1199 178 1203 183
rect 1 119 5 178
rect 1014 174 1066 178
rect 1199 176 1200 178
rect 1202 176 1203 178
rect 1102 171 1106 174
rect 1102 169 1103 171
rect 1105 169 1106 171
rect 1102 155 1106 169
rect 1199 155 1203 176
rect 1013 152 1017 155
rect 809 148 1017 152
rect 1063 151 1114 155
rect 306 145 311 148
rect 306 143 308 145
rect 310 143 311 145
rect 306 128 311 143
rect 556 144 561 145
rect 556 142 558 144
rect 560 142 561 144
rect 556 128 561 142
rect 809 128 813 148
rect 1063 128 1067 151
rect 1146 145 1150 147
rect 1146 143 1147 145
rect 1149 143 1150 145
rect 1146 135 1150 143
rect 1146 133 1147 135
rect 1149 133 1150 135
rect 1146 132 1150 133
rect 124 127 157 128
rect 124 125 125 127
rect 127 125 152 127
rect 154 125 157 127
rect 124 124 157 125
rect 181 127 220 128
rect 181 125 217 127
rect 219 125 220 127
rect 181 123 220 125
rect 279 127 312 128
rect 279 125 280 127
rect 282 125 307 127
rect 309 125 312 127
rect 279 124 312 125
rect 352 127 417 128
rect 352 125 353 127
rect 355 125 385 127
rect 387 125 412 127
rect 414 125 417 127
rect 352 124 417 125
rect 529 127 562 128
rect 529 125 530 127
rect 532 125 557 127
rect 559 125 562 127
rect 529 124 562 125
rect 602 127 667 128
rect 602 125 603 127
rect 605 125 635 127
rect 637 125 662 127
rect 664 125 667 127
rect 602 124 667 125
rect 779 127 813 128
rect 779 125 780 127
rect 782 125 807 127
rect 809 125 813 127
rect 779 124 813 125
rect 852 127 917 128
rect 852 125 853 127
rect 855 125 885 127
rect 887 125 912 127
rect 914 125 917 127
rect 852 124 917 125
rect 1029 127 1067 128
rect 1029 125 1030 127
rect 1032 125 1057 127
rect 1059 125 1067 127
rect 1029 124 1067 125
rect 1102 127 1167 128
rect 1102 125 1103 127
rect 1105 125 1135 127
rect 1137 125 1162 127
rect 1164 125 1167 127
rect 1102 124 1167 125
rect 181 120 186 123
rect 1 118 119 119
rect 1 116 116 118
rect 118 116 119 118
rect 1 115 119 116
rect 141 115 186 120
rect 1146 119 1150 120
rect 1146 117 1147 119
rect 1149 117 1150 119
rect 141 110 146 115
rect 141 108 143 110
rect 145 108 146 110
rect 141 107 146 108
rect 197 113 201 117
rect 197 111 198 113
rect 200 111 201 113
rect 84 101 105 103
rect 84 99 102 101
rect 104 99 105 101
rect 84 97 105 99
rect 84 75 89 97
rect 197 76 201 111
rect 1146 110 1150 117
rect 394 109 469 110
rect 394 107 395 109
rect 397 107 466 109
rect 468 107 469 109
rect 394 106 469 107
rect 646 109 719 110
rect 646 107 647 109
rect 649 107 716 109
rect 718 107 719 109
rect 646 106 719 107
rect 896 109 969 110
rect 896 107 897 109
rect 899 107 966 109
rect 968 107 969 109
rect 1146 108 1147 110
rect 1149 108 1150 110
rect 1146 107 1150 108
rect 896 106 969 107
rect 247 101 365 102
rect 247 99 248 101
rect 250 99 362 101
rect 364 99 365 101
rect 247 98 365 99
rect 457 101 461 102
rect 457 99 458 101
rect 460 99 461 101
rect 197 72 290 76
rect 457 75 461 99
rect 497 101 615 102
rect 497 99 498 101
rect 500 99 612 101
rect 614 99 615 101
rect 497 98 615 99
rect 707 101 711 102
rect 707 99 708 101
rect 710 99 711 101
rect 707 75 711 99
rect 747 101 865 102
rect 747 99 748 101
rect 750 99 862 101
rect 864 99 865 101
rect 747 98 865 99
rect 997 101 1115 102
rect 997 99 998 101
rect 1000 99 1112 101
rect 1114 99 1115 101
rect 997 98 1115 99
rect 39 55 157 56
rect 39 53 40 55
rect 42 53 154 55
rect 156 53 157 55
rect 39 52 157 53
rect 173 40 178 69
rect 286 56 290 72
rect 546 69 550 75
rect 530 65 550 69
rect 796 65 800 75
rect 286 55 407 56
rect 286 53 290 55
rect 292 53 404 55
rect 406 53 407 55
rect 286 52 407 53
rect 186 47 261 48
rect 186 45 187 47
rect 189 45 258 47
rect 260 45 261 47
rect 186 44 261 45
rect 104 38 178 40
rect 104 36 106 38
rect 108 36 178 38
rect 104 35 178 36
rect 286 40 290 52
rect 438 47 511 48
rect 438 45 439 47
rect 441 45 508 47
rect 510 45 511 47
rect 438 44 511 45
rect 530 40 534 65
rect 779 60 800 65
rect 539 55 657 56
rect 539 53 540 55
rect 542 53 654 55
rect 656 53 657 55
rect 539 52 657 53
rect 688 47 761 48
rect 688 45 689 47
rect 691 45 758 47
rect 760 45 761 47
rect 688 44 761 45
rect 779 40 784 60
rect 789 55 907 56
rect 789 53 790 55
rect 792 53 904 55
rect 906 53 907 55
rect 789 52 907 53
rect 938 46 942 47
rect 938 44 939 46
rect 941 44 942 46
rect 286 39 359 40
rect 286 37 356 39
rect 358 37 359 39
rect 286 35 359 37
rect 530 39 609 40
rect 530 37 606 39
rect 608 37 609 39
rect 530 36 609 37
rect 779 38 859 40
rect 779 36 856 38
rect 858 36 859 38
rect 779 34 859 36
rect 938 37 942 44
rect 938 35 939 37
rect 941 35 942 37
rect 938 34 942 35
rect 71 29 104 30
rect 71 27 72 29
rect 74 27 99 29
rect 101 27 104 29
rect 71 26 104 27
rect 144 29 209 30
rect 144 27 145 29
rect 147 27 177 29
rect 179 27 204 29
rect 206 27 209 29
rect 144 26 209 27
rect 321 29 354 30
rect 321 27 322 29
rect 324 27 349 29
rect 351 27 354 29
rect 321 26 354 27
rect 394 29 459 30
rect 394 27 395 29
rect 397 27 427 29
rect 429 27 454 29
rect 456 27 459 29
rect 394 26 459 27
rect 571 29 604 30
rect 571 27 572 29
rect 574 27 599 29
rect 601 27 604 29
rect 571 26 604 27
rect 644 29 709 30
rect 644 27 645 29
rect 647 27 677 29
rect 679 27 704 29
rect 706 27 709 29
rect 644 26 709 27
rect 821 29 854 30
rect 821 27 822 29
rect 824 27 849 29
rect 851 27 854 29
rect 821 26 854 27
rect 894 29 959 30
rect 894 27 895 29
rect 897 27 927 29
rect 929 27 954 29
rect 956 27 959 29
rect 894 26 959 27
rect 938 21 942 22
rect 938 19 939 21
rect 941 19 942 21
rect 938 11 942 19
rect 938 9 939 11
rect 941 9 942 11
rect 938 7 942 9
<< alu3 >>
rect 1102 190 1106 191
rect 1102 188 1103 190
rect 1105 188 1106 190
rect 1102 171 1106 188
rect 1102 169 1103 171
rect 1105 169 1106 171
rect 1102 168 1106 169
rect 1146 135 1150 136
rect 1146 133 1147 135
rect 1149 133 1150 135
rect 1146 119 1150 133
rect 1146 117 1147 119
rect 1149 117 1150 119
rect 1146 116 1150 117
rect 938 37 942 38
rect 938 35 939 37
rect 941 35 942 37
rect 938 21 942 35
rect 938 19 939 21
rect 941 19 942 21
rect 938 18 942 19
<< ptie >>
rect 43 413 49 415
rect 43 411 45 413
rect 47 411 49 413
rect 43 409 49 411
rect 83 413 89 415
rect 83 411 85 413
rect 87 411 89 413
rect 83 409 89 411
rect 154 413 160 415
rect 154 411 156 413
rect 158 411 160 413
rect 154 409 160 411
rect 195 413 201 415
rect 195 411 197 413
rect 199 411 201 413
rect 195 409 201 411
rect 525 415 531 417
rect 525 413 527 415
rect 529 413 531 415
rect 525 411 531 413
rect 565 415 571 417
rect 565 413 567 415
rect 569 413 571 415
rect 565 411 571 413
rect 636 415 642 417
rect 636 413 638 415
rect 640 413 642 415
rect 636 411 642 413
rect 677 415 683 417
rect 677 413 679 415
rect 681 413 683 415
rect 677 411 683 413
rect 730 415 736 417
rect 730 413 732 415
rect 734 413 736 415
rect 730 411 736 413
rect 770 415 776 417
rect 770 413 772 415
rect 774 413 776 415
rect 770 411 776 413
rect 841 415 847 417
rect 841 413 843 415
rect 845 413 847 415
rect 841 411 847 413
rect 882 415 888 417
rect 882 413 884 415
rect 886 413 888 415
rect 882 411 888 413
rect 15 281 21 283
rect 15 279 17 281
rect 19 279 21 281
rect 15 277 21 279
rect 83 281 89 283
rect 83 279 85 281
rect 87 279 89 281
rect 83 277 89 279
rect 95 281 101 283
rect 95 279 97 281
rect 99 279 101 281
rect 95 277 101 279
rect 136 281 142 283
rect 136 279 138 281
rect 140 279 142 281
rect 136 277 142 279
rect 497 283 503 285
rect 497 281 499 283
rect 501 281 503 283
rect 497 279 503 281
rect 565 283 571 285
rect 565 281 567 283
rect 569 281 571 283
rect 565 279 571 281
rect 577 283 583 285
rect 577 281 579 283
rect 581 281 583 283
rect 577 279 583 281
rect 618 283 624 285
rect 618 281 620 283
rect 622 281 624 283
rect 618 279 624 281
rect 702 283 708 285
rect 702 281 704 283
rect 706 281 708 283
rect 702 279 708 281
rect 770 283 776 285
rect 770 281 772 283
rect 774 281 776 283
rect 770 279 776 281
rect 782 283 788 285
rect 782 281 784 283
rect 786 281 788 283
rect 782 279 788 281
rect 823 283 829 285
rect 823 281 825 283
rect 827 281 829 283
rect 823 279 829 281
rect 1051 297 1057 299
rect 1051 295 1053 297
rect 1055 295 1057 297
rect 1051 293 1057 295
rect 1091 297 1097 299
rect 1091 295 1093 297
rect 1095 295 1097 297
rect 1091 293 1097 295
rect 1162 297 1168 299
rect 1162 295 1164 297
rect 1166 295 1168 297
rect 1162 293 1168 295
rect 1203 297 1209 299
rect 1203 295 1205 297
rect 1207 295 1209 297
rect 1203 293 1209 295
rect 2 165 8 167
rect 42 165 48 167
rect 2 163 4 165
rect 6 163 8 165
rect 2 161 8 163
rect 42 163 44 165
rect 46 163 48 165
rect 42 161 48 163
rect 83 165 89 167
rect 83 163 85 165
rect 87 163 89 165
rect 83 161 89 163
rect 147 165 153 167
rect 147 163 149 165
rect 151 163 153 165
rect 147 161 153 163
rect 188 165 194 167
rect 188 163 190 165
rect 192 163 194 165
rect 188 161 194 163
rect 252 165 258 167
rect 292 165 298 167
rect 252 163 254 165
rect 256 163 258 165
rect 252 161 258 163
rect 292 163 294 165
rect 296 163 298 165
rect 292 161 298 163
rect 333 165 339 167
rect 333 163 335 165
rect 337 163 339 165
rect 333 161 339 163
rect 397 165 403 167
rect 397 163 399 165
rect 401 163 403 165
rect 397 161 403 163
rect 438 165 444 167
rect 438 163 440 165
rect 442 163 444 165
rect 438 161 444 163
rect 502 165 508 167
rect 542 165 548 167
rect 502 163 504 165
rect 506 163 508 165
rect 502 161 508 163
rect 542 163 544 165
rect 546 163 548 165
rect 542 161 548 163
rect 583 165 589 167
rect 583 163 585 165
rect 587 163 589 165
rect 583 161 589 163
rect 647 165 653 167
rect 647 163 649 165
rect 651 163 653 165
rect 647 161 653 163
rect 688 165 694 167
rect 688 163 690 165
rect 692 163 694 165
rect 688 161 694 163
rect 752 165 758 167
rect 792 165 798 167
rect 752 163 754 165
rect 756 163 758 165
rect 752 161 758 163
rect 792 163 794 165
rect 796 163 798 165
rect 792 161 798 163
rect 833 165 839 167
rect 833 163 835 165
rect 837 163 839 165
rect 833 161 839 163
rect 897 165 903 167
rect 897 163 899 165
rect 901 163 903 165
rect 897 161 903 163
rect 938 165 944 167
rect 938 163 940 165
rect 942 163 944 165
rect 938 161 944 163
rect 1023 165 1029 167
rect 1023 163 1025 165
rect 1027 163 1029 165
rect 1023 161 1029 163
rect 1091 165 1097 167
rect 1091 163 1093 165
rect 1095 163 1097 165
rect 1091 161 1097 163
rect 1103 165 1109 167
rect 1103 163 1105 165
rect 1107 163 1109 165
rect 1103 161 1109 163
rect 1144 165 1150 167
rect 1144 163 1146 165
rect 1148 163 1150 165
rect 1144 161 1150 163
rect 101 144 107 146
rect 101 142 103 144
rect 105 142 107 144
rect 101 140 107 142
rect 142 144 148 146
rect 142 142 144 144
rect 146 142 148 144
rect 142 140 148 142
rect 216 144 222 146
rect 216 142 218 144
rect 220 142 222 144
rect 256 144 262 146
rect 256 142 258 144
rect 260 142 262 144
rect 216 140 222 142
rect 256 140 262 142
rect 297 144 303 146
rect 297 142 299 144
rect 301 142 303 144
rect 297 140 303 142
rect 361 144 367 146
rect 361 142 363 144
rect 365 142 367 144
rect 361 140 367 142
rect 402 144 408 146
rect 402 142 404 144
rect 406 142 408 144
rect 402 140 408 142
rect 466 144 472 146
rect 466 142 468 144
rect 470 142 472 144
rect 506 144 512 146
rect 506 142 508 144
rect 510 142 512 144
rect 466 140 472 142
rect 506 140 512 142
rect 547 144 553 146
rect 547 142 549 144
rect 551 142 553 144
rect 547 140 553 142
rect 611 144 617 146
rect 611 142 613 144
rect 615 142 617 144
rect 611 140 617 142
rect 652 144 658 146
rect 652 142 654 144
rect 656 142 658 144
rect 652 140 658 142
rect 716 144 722 146
rect 716 142 718 144
rect 720 142 722 144
rect 756 144 762 146
rect 756 142 758 144
rect 760 142 762 144
rect 716 140 722 142
rect 756 140 762 142
rect 797 144 803 146
rect 797 142 799 144
rect 801 142 803 144
rect 797 140 803 142
rect 861 144 867 146
rect 861 142 863 144
rect 865 142 867 144
rect 861 140 867 142
rect 902 144 908 146
rect 902 142 904 144
rect 906 142 908 144
rect 902 140 908 142
rect 966 144 972 146
rect 966 142 968 144
rect 970 142 972 144
rect 1006 144 1012 146
rect 1006 142 1008 144
rect 1010 142 1012 144
rect 966 140 972 142
rect 1006 140 1012 142
rect 1047 144 1053 146
rect 1047 142 1049 144
rect 1051 142 1053 144
rect 1047 140 1053 142
rect 1111 144 1117 146
rect 1111 142 1113 144
rect 1115 142 1117 144
rect 1111 140 1117 142
rect 1152 144 1158 146
rect 1152 142 1154 144
rect 1156 142 1158 144
rect 1152 140 1158 142
rect 8 12 14 14
rect 48 12 54 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 48 10 50 12
rect 52 10 54 12
rect 48 8 54 10
rect 89 12 95 14
rect 89 10 91 12
rect 93 10 95 12
rect 89 8 95 10
rect 153 12 159 14
rect 153 10 155 12
rect 157 10 159 12
rect 153 8 159 10
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
rect 258 12 264 14
rect 298 12 304 14
rect 258 10 260 12
rect 262 10 264 12
rect 258 8 264 10
rect 298 10 300 12
rect 302 10 304 12
rect 298 8 304 10
rect 339 12 345 14
rect 339 10 341 12
rect 343 10 345 12
rect 339 8 345 10
rect 403 12 409 14
rect 403 10 405 12
rect 407 10 409 12
rect 403 8 409 10
rect 444 12 450 14
rect 444 10 446 12
rect 448 10 450 12
rect 444 8 450 10
rect 508 12 514 14
rect 548 12 554 14
rect 508 10 510 12
rect 512 10 514 12
rect 508 8 514 10
rect 548 10 550 12
rect 552 10 554 12
rect 548 8 554 10
rect 589 12 595 14
rect 589 10 591 12
rect 593 10 595 12
rect 589 8 595 10
rect 653 12 659 14
rect 653 10 655 12
rect 657 10 659 12
rect 653 8 659 10
rect 694 12 700 14
rect 694 10 696 12
rect 698 10 700 12
rect 694 8 700 10
rect 758 12 764 14
rect 798 12 804 14
rect 758 10 760 12
rect 762 10 764 12
rect 758 8 764 10
rect 798 10 800 12
rect 802 10 804 12
rect 798 8 804 10
rect 839 12 845 14
rect 839 10 841 12
rect 843 10 845 12
rect 839 8 845 10
rect 903 12 909 14
rect 903 10 905 12
rect 907 10 909 12
rect 903 8 909 10
rect 944 12 950 14
rect 944 10 946 12
rect 948 10 950 12
rect 944 8 950 10
<< ntie >>
rect 43 353 49 355
rect 43 351 45 353
rect 47 351 49 353
rect 43 349 49 351
rect 83 353 89 355
rect 83 351 85 353
rect 87 351 89 353
rect 121 353 127 355
rect 83 349 89 351
rect 121 351 123 353
rect 125 351 127 353
rect 525 355 531 357
rect 195 353 201 355
rect 121 349 127 351
rect 195 351 197 353
rect 199 351 201 353
rect 525 353 527 355
rect 529 353 531 355
rect 525 351 531 353
rect 565 355 571 357
rect 565 353 567 355
rect 569 353 571 355
rect 603 355 609 357
rect 565 351 571 353
rect 195 349 201 351
rect 603 353 605 355
rect 607 353 609 355
rect 677 355 683 357
rect 603 351 609 353
rect 677 353 679 355
rect 681 353 683 355
rect 677 351 683 353
rect 730 355 736 357
rect 730 353 732 355
rect 734 353 736 355
rect 730 351 736 353
rect 770 355 776 357
rect 770 353 772 355
rect 774 353 776 355
rect 808 355 814 357
rect 770 351 776 353
rect 808 353 810 355
rect 812 353 814 355
rect 882 355 888 357
rect 808 351 814 353
rect 882 353 884 355
rect 886 353 888 355
rect 882 351 888 353
rect 15 341 21 343
rect 15 339 17 341
rect 19 339 21 341
rect 15 337 21 339
rect 83 341 89 343
rect 83 339 85 341
rect 87 339 89 341
rect 83 337 89 339
rect 95 341 101 343
rect 95 339 97 341
rect 99 339 101 341
rect 169 341 175 343
rect 95 337 101 339
rect 169 339 171 341
rect 173 339 175 341
rect 497 343 503 345
rect 497 341 499 343
rect 501 341 503 343
rect 169 337 175 339
rect 497 339 503 341
rect 565 343 571 345
rect 565 341 567 343
rect 569 341 571 343
rect 565 339 571 341
rect 577 343 583 345
rect 577 341 579 343
rect 581 341 583 343
rect 651 343 657 345
rect 577 339 583 341
rect 651 341 653 343
rect 655 341 657 343
rect 702 343 708 345
rect 651 339 657 341
rect 702 341 704 343
rect 706 341 708 343
rect 702 339 708 341
rect 770 343 776 345
rect 770 341 772 343
rect 774 341 776 343
rect 770 339 776 341
rect 782 343 788 345
rect 782 341 784 343
rect 786 341 788 343
rect 856 343 862 345
rect 782 339 788 341
rect 856 341 858 343
rect 860 341 862 343
rect 856 339 862 341
rect 1051 237 1057 239
rect 1051 235 1053 237
rect 1055 235 1057 237
rect 1051 233 1057 235
rect 1091 237 1097 239
rect 1091 235 1093 237
rect 1095 235 1097 237
rect 1129 237 1135 239
rect 1091 233 1097 235
rect 1129 235 1131 237
rect 1133 235 1135 237
rect 1203 237 1209 239
rect 1129 233 1135 235
rect 1203 235 1205 237
rect 1207 235 1209 237
rect 1203 233 1209 235
rect 2 225 8 227
rect 2 223 4 225
rect 6 223 8 225
rect 42 225 48 227
rect 2 221 8 223
rect 42 223 44 225
rect 46 223 48 225
rect 116 225 122 227
rect 42 221 48 223
rect 116 223 118 225
rect 120 223 122 225
rect 147 225 153 227
rect 116 221 122 223
rect 147 223 149 225
rect 151 223 153 225
rect 221 225 227 227
rect 147 221 153 223
rect 221 223 223 225
rect 225 223 227 225
rect 252 225 258 227
rect 221 221 227 223
rect 252 223 254 225
rect 256 223 258 225
rect 292 225 298 227
rect 252 221 258 223
rect 292 223 294 225
rect 296 223 298 225
rect 366 225 372 227
rect 292 221 298 223
rect 366 223 368 225
rect 370 223 372 225
rect 397 225 403 227
rect 366 221 372 223
rect 397 223 399 225
rect 401 223 403 225
rect 471 225 477 227
rect 397 221 403 223
rect 471 223 473 225
rect 475 223 477 225
rect 502 225 508 227
rect 471 221 477 223
rect 502 223 504 225
rect 506 223 508 225
rect 542 225 548 227
rect 502 221 508 223
rect 542 223 544 225
rect 546 223 548 225
rect 616 225 622 227
rect 542 221 548 223
rect 616 223 618 225
rect 620 223 622 225
rect 647 225 653 227
rect 616 221 622 223
rect 647 223 649 225
rect 651 223 653 225
rect 721 225 727 227
rect 647 221 653 223
rect 721 223 723 225
rect 725 223 727 225
rect 752 225 758 227
rect 721 221 727 223
rect 752 223 754 225
rect 756 223 758 225
rect 792 225 798 227
rect 752 221 758 223
rect 792 223 794 225
rect 796 223 798 225
rect 866 225 872 227
rect 792 221 798 223
rect 866 223 868 225
rect 870 223 872 225
rect 897 225 903 227
rect 866 221 872 223
rect 897 223 899 225
rect 901 223 903 225
rect 971 225 977 227
rect 897 221 903 223
rect 971 223 973 225
rect 975 223 977 225
rect 1023 225 1029 227
rect 971 221 977 223
rect 1023 223 1025 225
rect 1027 223 1029 225
rect 1023 221 1029 223
rect 1091 225 1097 227
rect 1091 223 1093 225
rect 1095 223 1097 225
rect 1091 221 1097 223
rect 1103 225 1109 227
rect 1103 223 1105 225
rect 1107 223 1109 225
rect 1177 225 1183 227
rect 1103 221 1109 223
rect 1177 223 1179 225
rect 1181 223 1183 225
rect 1177 221 1183 223
rect 101 84 107 86
rect 101 82 103 84
rect 105 82 107 84
rect 175 84 181 86
rect 101 80 107 82
rect 175 82 177 84
rect 179 82 181 84
rect 216 84 222 86
rect 175 80 181 82
rect 216 82 218 84
rect 220 82 222 84
rect 256 84 262 86
rect 216 80 222 82
rect 256 82 258 84
rect 260 82 262 84
rect 330 84 336 86
rect 256 80 262 82
rect 330 82 332 84
rect 334 82 336 84
rect 361 84 367 86
rect 330 80 336 82
rect 361 82 363 84
rect 365 82 367 84
rect 435 84 441 86
rect 361 80 367 82
rect 435 82 437 84
rect 439 82 441 84
rect 466 84 472 86
rect 435 80 441 82
rect 466 82 468 84
rect 470 82 472 84
rect 506 84 512 86
rect 466 80 472 82
rect 506 82 508 84
rect 510 82 512 84
rect 580 84 586 86
rect 506 80 512 82
rect 580 82 582 84
rect 584 82 586 84
rect 611 84 617 86
rect 580 80 586 82
rect 611 82 613 84
rect 615 82 617 84
rect 685 84 691 86
rect 611 80 617 82
rect 685 82 687 84
rect 689 82 691 84
rect 716 84 722 86
rect 685 80 691 82
rect 716 82 718 84
rect 720 82 722 84
rect 756 84 762 86
rect 716 80 722 82
rect 756 82 758 84
rect 760 82 762 84
rect 830 84 836 86
rect 756 80 762 82
rect 830 82 832 84
rect 834 82 836 84
rect 861 84 867 86
rect 830 80 836 82
rect 861 82 863 84
rect 865 82 867 84
rect 935 84 941 86
rect 861 80 867 82
rect 935 82 937 84
rect 939 82 941 84
rect 966 84 972 86
rect 935 80 941 82
rect 966 82 968 84
rect 970 82 972 84
rect 1006 84 1012 86
rect 966 80 972 82
rect 1006 82 1008 84
rect 1010 82 1012 84
rect 1080 84 1086 86
rect 1006 80 1012 82
rect 1080 82 1082 84
rect 1084 82 1086 84
rect 1111 84 1117 86
rect 1080 80 1086 82
rect 1111 82 1113 84
rect 1115 82 1117 84
rect 1185 84 1191 86
rect 1111 80 1117 82
rect 1185 82 1187 84
rect 1189 82 1191 84
rect 1185 80 1191 82
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 48 72 54 74
rect 8 68 14 70
rect 48 70 50 72
rect 52 70 54 72
rect 122 72 128 74
rect 48 68 54 70
rect 122 70 124 72
rect 126 70 128 72
rect 153 72 159 74
rect 122 68 128 70
rect 153 70 155 72
rect 157 70 159 72
rect 227 72 233 74
rect 153 68 159 70
rect 227 70 229 72
rect 231 70 233 72
rect 258 72 264 74
rect 227 68 233 70
rect 258 70 260 72
rect 262 70 264 72
rect 298 72 304 74
rect 258 68 264 70
rect 298 70 300 72
rect 302 70 304 72
rect 372 72 378 74
rect 298 68 304 70
rect 372 70 374 72
rect 376 70 378 72
rect 403 72 409 74
rect 372 68 378 70
rect 403 70 405 72
rect 407 70 409 72
rect 477 72 483 74
rect 403 68 409 70
rect 477 70 479 72
rect 481 70 483 72
rect 508 72 514 74
rect 477 68 483 70
rect 508 70 510 72
rect 512 70 514 72
rect 548 72 554 74
rect 508 68 514 70
rect 548 70 550 72
rect 552 70 554 72
rect 622 72 628 74
rect 548 68 554 70
rect 622 70 624 72
rect 626 70 628 72
rect 653 72 659 74
rect 622 68 628 70
rect 653 70 655 72
rect 657 70 659 72
rect 727 72 733 74
rect 653 68 659 70
rect 727 70 729 72
rect 731 70 733 72
rect 758 72 764 74
rect 727 68 733 70
rect 758 70 760 72
rect 762 70 764 72
rect 798 72 804 74
rect 758 68 764 70
rect 798 70 800 72
rect 802 70 804 72
rect 872 72 878 74
rect 798 68 804 70
rect 872 70 874 72
rect 876 70 878 72
rect 903 72 909 74
rect 872 68 878 70
rect 903 70 905 72
rect 907 70 909 72
rect 977 72 983 74
rect 903 68 909 70
rect 977 70 979 72
rect 981 70 983 72
rect 977 68 983 70
<< nmos >>
rect 21 394 23 405
rect 28 394 30 405
rect 41 394 43 403
rect 61 394 63 405
rect 68 394 70 405
rect 81 394 83 403
rect 109 397 111 409
rect 116 397 118 409
rect 126 397 128 406
rect 136 397 138 406
rect 152 392 154 401
rect 173 394 175 405
rect 180 394 182 405
rect 193 394 195 403
rect 503 396 505 407
rect 510 396 512 407
rect 523 396 525 405
rect 543 396 545 407
rect 550 396 552 407
rect 563 396 565 405
rect 591 399 593 411
rect 598 399 600 411
rect 608 399 610 408
rect 618 399 620 408
rect 634 394 636 403
rect 655 396 657 407
rect 662 396 664 407
rect 675 396 677 405
rect 708 396 710 407
rect 715 396 717 407
rect 728 396 730 405
rect 748 396 750 407
rect 755 396 757 407
rect 768 396 770 405
rect 796 399 798 411
rect 803 399 805 411
rect 813 399 815 408
rect 823 399 825 408
rect 839 394 841 403
rect 860 396 862 407
rect 867 396 869 407
rect 880 396 882 405
rect 21 289 23 298
rect 34 287 36 298
rect 41 287 43 298
rect 61 287 63 298
rect 68 287 70 298
rect 81 289 83 298
rect 101 289 103 298
rect 114 287 116 298
rect 121 287 123 298
rect 142 291 144 300
rect 158 286 160 295
rect 168 286 170 295
rect 178 283 180 295
rect 185 283 187 295
rect 503 291 505 300
rect 516 289 518 300
rect 523 289 525 300
rect 543 289 545 300
rect 550 289 552 300
rect 563 291 565 300
rect 583 291 585 300
rect 596 289 598 300
rect 603 289 605 300
rect 624 293 626 302
rect 640 288 642 297
rect 650 288 652 297
rect 660 285 662 297
rect 667 285 669 297
rect 708 291 710 300
rect 721 289 723 300
rect 728 289 730 300
rect 748 289 750 300
rect 755 289 757 300
rect 768 291 770 300
rect 788 291 790 300
rect 801 289 803 300
rect 808 289 810 300
rect 829 293 831 302
rect 845 288 847 297
rect 855 288 857 297
rect 865 285 867 297
rect 872 285 874 297
rect 1029 278 1031 289
rect 1036 278 1038 289
rect 1049 278 1051 287
rect 1069 278 1071 289
rect 1076 278 1078 289
rect 1089 278 1091 287
rect 1117 281 1119 293
rect 1124 281 1126 293
rect 1134 281 1136 290
rect 1144 281 1146 290
rect 1160 276 1162 285
rect 1181 278 1183 289
rect 1188 278 1190 289
rect 1201 278 1203 287
rect 8 175 10 184
rect 18 178 20 184
rect 28 178 30 184
rect 48 173 50 182
rect 61 171 63 182
rect 68 171 70 182
rect 89 175 91 184
rect 105 170 107 179
rect 115 170 117 179
rect 125 167 127 179
rect 132 167 134 179
rect 153 173 155 182
rect 166 171 168 182
rect 173 171 175 182
rect 194 175 196 184
rect 210 170 212 179
rect 220 170 222 179
rect 230 167 232 179
rect 237 167 239 179
rect 258 175 260 184
rect 268 178 270 184
rect 278 178 280 184
rect 298 173 300 182
rect 311 171 313 182
rect 318 171 320 182
rect 339 175 341 184
rect 355 170 357 179
rect 365 170 367 179
rect 375 167 377 179
rect 382 167 384 179
rect 403 173 405 182
rect 416 171 418 182
rect 423 171 425 182
rect 444 175 446 184
rect 460 170 462 179
rect 470 170 472 179
rect 480 167 482 179
rect 487 167 489 179
rect 508 175 510 184
rect 518 178 520 184
rect 528 178 530 184
rect 548 173 550 182
rect 561 171 563 182
rect 568 171 570 182
rect 589 175 591 184
rect 605 170 607 179
rect 615 170 617 179
rect 625 167 627 179
rect 632 167 634 179
rect 653 173 655 182
rect 666 171 668 182
rect 673 171 675 182
rect 694 175 696 184
rect 710 170 712 179
rect 720 170 722 179
rect 730 167 732 179
rect 737 167 739 179
rect 758 175 760 184
rect 768 178 770 184
rect 778 178 780 184
rect 798 173 800 182
rect 811 171 813 182
rect 818 171 820 182
rect 839 175 841 184
rect 855 170 857 179
rect 865 170 867 179
rect 875 167 877 179
rect 882 167 884 179
rect 903 173 905 182
rect 916 171 918 182
rect 923 171 925 182
rect 944 175 946 184
rect 960 170 962 179
rect 970 170 972 179
rect 980 167 982 179
rect 987 167 989 179
rect 1029 173 1031 182
rect 1042 171 1044 182
rect 1049 171 1051 182
rect 1069 171 1071 182
rect 1076 171 1078 182
rect 1089 173 1091 182
rect 1109 173 1111 182
rect 1122 171 1124 182
rect 1129 171 1131 182
rect 1150 175 1152 184
rect 1166 170 1168 179
rect 1176 170 1178 179
rect 1186 167 1188 179
rect 1193 167 1195 179
rect 107 125 109 134
rect 120 125 122 136
rect 127 125 129 136
rect 148 123 150 132
rect 164 128 166 137
rect 174 128 176 137
rect 184 128 186 140
rect 191 128 193 140
rect 222 123 224 132
rect 232 123 234 129
rect 242 123 244 129
rect 262 125 264 134
rect 275 125 277 136
rect 282 125 284 136
rect 303 123 305 132
rect 319 128 321 137
rect 329 128 331 137
rect 339 128 341 140
rect 346 128 348 140
rect 367 125 369 134
rect 380 125 382 136
rect 387 125 389 136
rect 408 123 410 132
rect 424 128 426 137
rect 434 128 436 137
rect 444 128 446 140
rect 451 128 453 140
rect 472 123 474 132
rect 482 123 484 129
rect 492 123 494 129
rect 512 125 514 134
rect 525 125 527 136
rect 532 125 534 136
rect 553 123 555 132
rect 569 128 571 137
rect 579 128 581 137
rect 589 128 591 140
rect 596 128 598 140
rect 617 125 619 134
rect 630 125 632 136
rect 637 125 639 136
rect 658 123 660 132
rect 674 128 676 137
rect 684 128 686 137
rect 694 128 696 140
rect 701 128 703 140
rect 722 123 724 132
rect 732 123 734 129
rect 742 123 744 129
rect 762 125 764 134
rect 775 125 777 136
rect 782 125 784 136
rect 803 123 805 132
rect 819 128 821 137
rect 829 128 831 137
rect 839 128 841 140
rect 846 128 848 140
rect 867 125 869 134
rect 880 125 882 136
rect 887 125 889 136
rect 908 123 910 132
rect 924 128 926 137
rect 934 128 936 137
rect 944 128 946 140
rect 951 128 953 140
rect 972 123 974 132
rect 982 123 984 129
rect 992 123 994 129
rect 1012 125 1014 134
rect 1025 125 1027 136
rect 1032 125 1034 136
rect 1053 123 1055 132
rect 1069 128 1071 137
rect 1079 128 1081 137
rect 1089 128 1091 140
rect 1096 128 1098 140
rect 1117 125 1119 134
rect 1130 125 1132 136
rect 1137 125 1139 136
rect 1158 123 1160 132
rect 1174 128 1176 137
rect 1184 128 1186 137
rect 1194 128 1196 140
rect 1201 128 1203 140
rect 14 22 16 31
rect 24 25 26 31
rect 34 25 36 31
rect 54 20 56 29
rect 67 18 69 29
rect 74 18 76 29
rect 95 22 97 31
rect 111 17 113 26
rect 121 17 123 26
rect 131 14 133 26
rect 138 14 140 26
rect 159 20 161 29
rect 172 18 174 29
rect 179 18 181 29
rect 200 22 202 31
rect 216 17 218 26
rect 226 17 228 26
rect 236 14 238 26
rect 243 14 245 26
rect 264 22 266 31
rect 274 25 276 31
rect 284 25 286 31
rect 304 20 306 29
rect 317 18 319 29
rect 324 18 326 29
rect 345 22 347 31
rect 361 17 363 26
rect 371 17 373 26
rect 381 14 383 26
rect 388 14 390 26
rect 409 20 411 29
rect 422 18 424 29
rect 429 18 431 29
rect 450 22 452 31
rect 466 17 468 26
rect 476 17 478 26
rect 486 14 488 26
rect 493 14 495 26
rect 514 22 516 31
rect 524 25 526 31
rect 534 25 536 31
rect 554 20 556 29
rect 567 18 569 29
rect 574 18 576 29
rect 595 22 597 31
rect 611 17 613 26
rect 621 17 623 26
rect 631 14 633 26
rect 638 14 640 26
rect 659 20 661 29
rect 672 18 674 29
rect 679 18 681 29
rect 700 22 702 31
rect 716 17 718 26
rect 726 17 728 26
rect 736 14 738 26
rect 743 14 745 26
rect 764 22 766 31
rect 774 25 776 31
rect 784 25 786 31
rect 804 20 806 29
rect 817 18 819 29
rect 824 18 826 29
rect 845 22 847 31
rect 861 17 863 26
rect 871 17 873 26
rect 881 14 883 26
rect 888 14 890 26
rect 909 20 911 29
rect 922 18 924 29
rect 929 18 931 29
rect 950 22 952 31
rect 966 17 968 26
rect 976 17 978 26
rect 986 14 988 26
rect 993 14 995 26
<< pmos >>
rect 21 359 23 372
rect 31 359 33 372
rect 41 361 43 379
rect 61 359 63 372
rect 71 359 73 372
rect 81 361 83 379
rect 108 352 110 379
rect 118 361 120 379
rect 128 361 130 379
rect 144 352 146 379
rect 173 359 175 372
rect 183 359 185 372
rect 193 361 195 379
rect 503 361 505 374
rect 513 361 515 374
rect 523 363 525 381
rect 543 361 545 374
rect 553 361 555 374
rect 563 363 565 381
rect 590 354 592 381
rect 600 363 602 381
rect 610 363 612 381
rect 626 354 628 381
rect 655 361 657 374
rect 665 361 667 374
rect 675 363 677 381
rect 708 361 710 374
rect 718 361 720 374
rect 728 363 730 381
rect 748 361 750 374
rect 758 361 760 374
rect 768 363 770 381
rect 795 354 797 381
rect 805 363 807 381
rect 815 363 817 381
rect 831 354 833 381
rect 860 361 862 374
rect 870 361 872 374
rect 880 363 882 381
rect 21 313 23 331
rect 31 320 33 333
rect 41 320 43 333
rect 61 320 63 333
rect 71 320 73 333
rect 81 313 83 331
rect 101 313 103 331
rect 111 320 113 333
rect 121 320 123 333
rect 150 313 152 340
rect 166 313 168 331
rect 176 313 178 331
rect 186 313 188 340
rect 503 315 505 333
rect 513 322 515 335
rect 523 322 525 335
rect 543 322 545 335
rect 553 322 555 335
rect 563 315 565 333
rect 583 315 585 333
rect 593 322 595 335
rect 603 322 605 335
rect 632 315 634 342
rect 648 315 650 333
rect 658 315 660 333
rect 668 315 670 342
rect 708 315 710 333
rect 718 322 720 335
rect 728 322 730 335
rect 748 322 750 335
rect 758 322 760 335
rect 768 315 770 333
rect 788 315 790 333
rect 798 322 800 335
rect 808 322 810 335
rect 837 315 839 342
rect 853 315 855 333
rect 863 315 865 333
rect 873 315 875 342
rect 1029 243 1031 256
rect 1039 243 1041 256
rect 1049 245 1051 263
rect 1069 243 1071 256
rect 1079 243 1081 256
rect 1089 245 1091 263
rect 1116 236 1118 263
rect 1126 245 1128 263
rect 1136 245 1138 263
rect 1152 236 1154 263
rect 1181 243 1183 256
rect 1191 243 1193 256
rect 1201 245 1203 263
rect 8 196 10 214
rect 21 203 23 224
rect 28 203 30 224
rect 48 197 50 215
rect 58 204 60 217
rect 68 204 70 217
rect 97 197 99 224
rect 113 197 115 215
rect 123 197 125 215
rect 133 197 135 224
rect 153 197 155 215
rect 163 204 165 217
rect 173 204 175 217
rect 202 197 204 224
rect 218 197 220 215
rect 228 197 230 215
rect 238 197 240 224
rect 258 196 260 214
rect 271 203 273 224
rect 278 203 280 224
rect 298 197 300 215
rect 308 204 310 217
rect 318 204 320 217
rect 347 197 349 224
rect 363 197 365 215
rect 373 197 375 215
rect 383 197 385 224
rect 403 197 405 215
rect 413 204 415 217
rect 423 204 425 217
rect 452 197 454 224
rect 468 197 470 215
rect 478 197 480 215
rect 488 197 490 224
rect 508 196 510 214
rect 521 203 523 224
rect 528 203 530 224
rect 548 197 550 215
rect 558 204 560 217
rect 568 204 570 217
rect 597 197 599 224
rect 613 197 615 215
rect 623 197 625 215
rect 633 197 635 224
rect 653 197 655 215
rect 663 204 665 217
rect 673 204 675 217
rect 702 197 704 224
rect 718 197 720 215
rect 728 197 730 215
rect 738 197 740 224
rect 758 196 760 214
rect 771 203 773 224
rect 778 203 780 224
rect 798 197 800 215
rect 808 204 810 217
rect 818 204 820 217
rect 847 197 849 224
rect 863 197 865 215
rect 873 197 875 215
rect 883 197 885 224
rect 903 197 905 215
rect 913 204 915 217
rect 923 204 925 217
rect 952 197 954 224
rect 968 197 970 215
rect 978 197 980 215
rect 988 197 990 224
rect 1029 197 1031 215
rect 1039 204 1041 217
rect 1049 204 1051 217
rect 1069 204 1071 217
rect 1079 204 1081 217
rect 1089 197 1091 215
rect 1109 197 1111 215
rect 1119 204 1121 217
rect 1129 204 1131 217
rect 1158 197 1160 224
rect 1174 197 1176 215
rect 1184 197 1186 215
rect 1194 197 1196 224
rect 107 92 109 110
rect 117 90 119 103
rect 127 90 129 103
rect 156 83 158 110
rect 172 92 174 110
rect 182 92 184 110
rect 192 83 194 110
rect 222 93 224 111
rect 235 83 237 104
rect 242 83 244 104
rect 262 92 264 110
rect 272 90 274 103
rect 282 90 284 103
rect 311 83 313 110
rect 327 92 329 110
rect 337 92 339 110
rect 347 83 349 110
rect 367 92 369 110
rect 377 90 379 103
rect 387 90 389 103
rect 416 83 418 110
rect 432 92 434 110
rect 442 92 444 110
rect 452 83 454 110
rect 472 93 474 111
rect 485 83 487 104
rect 492 83 494 104
rect 512 92 514 110
rect 522 90 524 103
rect 532 90 534 103
rect 561 83 563 110
rect 577 92 579 110
rect 587 92 589 110
rect 597 83 599 110
rect 617 92 619 110
rect 627 90 629 103
rect 637 90 639 103
rect 666 83 668 110
rect 682 92 684 110
rect 692 92 694 110
rect 702 83 704 110
rect 722 93 724 111
rect 735 83 737 104
rect 742 83 744 104
rect 762 92 764 110
rect 772 90 774 103
rect 782 90 784 103
rect 811 83 813 110
rect 827 92 829 110
rect 837 92 839 110
rect 847 83 849 110
rect 867 92 869 110
rect 877 90 879 103
rect 887 90 889 103
rect 916 83 918 110
rect 932 92 934 110
rect 942 92 944 110
rect 952 83 954 110
rect 972 93 974 111
rect 985 83 987 104
rect 992 83 994 104
rect 1012 92 1014 110
rect 1022 90 1024 103
rect 1032 90 1034 103
rect 1061 83 1063 110
rect 1077 92 1079 110
rect 1087 92 1089 110
rect 1097 83 1099 110
rect 1117 92 1119 110
rect 1127 90 1129 103
rect 1137 90 1139 103
rect 1166 83 1168 110
rect 1182 92 1184 110
rect 1192 92 1194 110
rect 1202 83 1204 110
rect 14 43 16 61
rect 27 50 29 71
rect 34 50 36 71
rect 54 44 56 62
rect 64 51 66 64
rect 74 51 76 64
rect 103 44 105 71
rect 119 44 121 62
rect 129 44 131 62
rect 139 44 141 71
rect 159 44 161 62
rect 169 51 171 64
rect 179 51 181 64
rect 208 44 210 71
rect 224 44 226 62
rect 234 44 236 62
rect 244 44 246 71
rect 264 43 266 61
rect 277 50 279 71
rect 284 50 286 71
rect 304 44 306 62
rect 314 51 316 64
rect 324 51 326 64
rect 353 44 355 71
rect 369 44 371 62
rect 379 44 381 62
rect 389 44 391 71
rect 409 44 411 62
rect 419 51 421 64
rect 429 51 431 64
rect 458 44 460 71
rect 474 44 476 62
rect 484 44 486 62
rect 494 44 496 71
rect 514 43 516 61
rect 527 50 529 71
rect 534 50 536 71
rect 554 44 556 62
rect 564 51 566 64
rect 574 51 576 64
rect 603 44 605 71
rect 619 44 621 62
rect 629 44 631 62
rect 639 44 641 71
rect 659 44 661 62
rect 669 51 671 64
rect 679 51 681 64
rect 708 44 710 71
rect 724 44 726 62
rect 734 44 736 62
rect 744 44 746 71
rect 764 43 766 61
rect 777 50 779 71
rect 784 50 786 71
rect 804 44 806 62
rect 814 51 816 64
rect 824 51 826 64
rect 853 44 855 71
rect 869 44 871 62
rect 879 44 881 62
rect 889 44 891 71
rect 909 44 911 62
rect 919 51 921 64
rect 929 51 931 64
rect 958 44 960 71
rect 974 44 976 62
rect 984 44 986 62
rect 994 44 996 71
<< polyct0 >>
rect 39 385 41 387
rect 79 385 81 387
rect 110 384 112 386
rect 120 385 122 387
rect 191 385 193 387
rect 521 387 523 389
rect 561 387 563 389
rect 592 386 594 388
rect 602 387 604 389
rect 673 387 675 389
rect 726 387 728 389
rect 766 387 768 389
rect 797 386 799 388
rect 807 387 809 389
rect 878 387 880 389
rect 23 305 25 307
rect 79 305 81 307
rect 103 305 105 307
rect 174 305 176 307
rect 184 306 186 308
rect 505 307 507 309
rect 561 307 563 309
rect 585 307 587 309
rect 656 307 658 309
rect 666 308 668 310
rect 710 307 712 309
rect 766 307 768 309
rect 790 307 792 309
rect 861 307 863 309
rect 871 308 873 310
rect 1047 269 1049 271
rect 1087 269 1089 271
rect 1118 268 1120 270
rect 1128 269 1130 271
rect 1199 269 1201 271
rect 10 189 12 191
rect 50 189 52 191
rect 121 189 123 191
rect 131 190 133 192
rect 155 189 157 191
rect 226 189 228 191
rect 236 190 238 192
rect 260 189 262 191
rect 300 189 302 191
rect 371 189 373 191
rect 381 190 383 192
rect 405 189 407 191
rect 476 189 478 191
rect 486 190 488 192
rect 510 189 512 191
rect 550 189 552 191
rect 621 189 623 191
rect 631 190 633 192
rect 655 189 657 191
rect 726 189 728 191
rect 736 190 738 192
rect 760 189 762 191
rect 800 189 802 191
rect 871 189 873 191
rect 881 190 883 192
rect 905 189 907 191
rect 976 189 978 191
rect 986 190 988 192
rect 1031 189 1033 191
rect 1087 189 1089 191
rect 1111 189 1113 191
rect 1182 189 1184 191
rect 1192 190 1194 192
rect 109 116 111 118
rect 180 116 182 118
rect 190 115 192 117
rect 224 116 226 118
rect 264 116 266 118
rect 335 116 337 118
rect 345 115 347 117
rect 369 116 371 118
rect 440 116 442 118
rect 450 115 452 117
rect 474 116 476 118
rect 514 116 516 118
rect 585 116 587 118
rect 595 115 597 117
rect 619 116 621 118
rect 690 116 692 118
rect 700 115 702 117
rect 724 116 726 118
rect 764 116 766 118
rect 835 116 837 118
rect 845 115 847 117
rect 869 116 871 118
rect 940 116 942 118
rect 950 115 952 117
rect 974 116 976 118
rect 1014 116 1016 118
rect 1085 116 1087 118
rect 1095 115 1097 117
rect 1119 116 1121 118
rect 1190 116 1192 118
rect 1200 115 1202 117
rect 16 36 18 38
rect 56 36 58 38
rect 127 36 129 38
rect 137 37 139 39
rect 161 36 163 38
rect 232 36 234 38
rect 242 37 244 39
rect 266 36 268 38
rect 306 36 308 38
rect 377 36 379 38
rect 387 37 389 39
rect 411 36 413 38
rect 482 36 484 38
rect 492 37 494 39
rect 516 36 518 38
rect 556 36 558 38
rect 627 36 629 38
rect 637 37 639 39
rect 661 36 663 38
rect 732 36 734 38
rect 742 37 744 39
rect 766 36 768 38
rect 806 36 808 38
rect 877 36 879 38
rect 887 37 889 39
rect 911 36 913 38
rect 982 36 984 38
rect 992 37 994 39
<< polyct1 >>
rect 29 385 31 387
rect 19 377 21 379
rect 69 385 71 387
rect 141 390 143 392
rect 59 377 61 379
rect 181 385 183 387
rect 511 387 513 389
rect 157 377 159 379
rect 171 377 173 379
rect 501 379 503 381
rect 551 387 553 389
rect 623 392 625 394
rect 541 379 543 381
rect 663 387 665 389
rect 639 379 641 381
rect 653 379 655 381
rect 716 387 718 389
rect 706 379 708 381
rect 756 387 758 389
rect 828 392 830 394
rect 746 379 748 381
rect 868 387 870 389
rect 844 379 846 381
rect 858 379 860 381
rect 43 313 45 315
rect 59 313 61 315
rect 33 305 35 307
rect 69 305 71 307
rect 123 313 125 315
rect 137 313 139 315
rect 113 305 115 307
rect 525 315 527 317
rect 541 315 543 317
rect 515 307 517 309
rect 153 300 155 302
rect 551 307 553 309
rect 605 315 607 317
rect 619 315 621 317
rect 595 307 597 309
rect 730 315 732 317
rect 746 315 748 317
rect 635 302 637 304
rect 720 307 722 309
rect 756 307 758 309
rect 810 315 812 317
rect 824 315 826 317
rect 800 307 802 309
rect 840 302 842 304
rect 1037 269 1039 271
rect 1027 261 1029 263
rect 1077 269 1079 271
rect 1149 274 1151 276
rect 1067 261 1069 263
rect 1189 269 1191 271
rect 1165 261 1167 263
rect 1179 261 1181 263
rect 30 196 32 198
rect 20 189 22 191
rect 70 197 72 199
rect 84 197 86 199
rect 60 189 62 191
rect 175 197 177 199
rect 189 197 191 199
rect 100 184 102 186
rect 165 189 167 191
rect 280 196 282 198
rect 205 184 207 186
rect 270 189 272 191
rect 320 197 322 199
rect 334 197 336 199
rect 310 189 312 191
rect 425 197 427 199
rect 439 197 441 199
rect 350 184 352 186
rect 415 189 417 191
rect 530 196 532 198
rect 455 184 457 186
rect 520 189 522 191
rect 570 197 572 199
rect 584 197 586 199
rect 560 189 562 191
rect 675 197 677 199
rect 689 197 691 199
rect 600 184 602 186
rect 665 189 667 191
rect 780 196 782 198
rect 705 184 707 186
rect 770 189 772 191
rect 820 197 822 199
rect 834 197 836 199
rect 810 189 812 191
rect 925 197 927 199
rect 939 197 941 199
rect 850 184 852 186
rect 915 189 917 191
rect 1051 197 1053 199
rect 1067 197 1069 199
rect 955 184 957 186
rect 1041 189 1043 191
rect 1077 189 1079 191
rect 1131 197 1133 199
rect 1145 197 1147 199
rect 1121 189 1123 191
rect 1161 184 1163 186
rect 119 116 121 118
rect 159 121 161 123
rect 129 108 131 110
rect 234 116 236 118
rect 143 108 145 110
rect 274 116 276 118
rect 244 109 246 111
rect 314 121 316 123
rect 284 108 286 110
rect 379 116 381 118
rect 298 108 300 110
rect 419 121 421 123
rect 389 108 391 110
rect 484 116 486 118
rect 403 108 405 110
rect 524 116 526 118
rect 494 109 496 111
rect 564 121 566 123
rect 534 108 536 110
rect 629 116 631 118
rect 548 108 550 110
rect 669 121 671 123
rect 639 108 641 110
rect 734 116 736 118
rect 653 108 655 110
rect 774 116 776 118
rect 744 109 746 111
rect 814 121 816 123
rect 784 108 786 110
rect 879 116 881 118
rect 798 108 800 110
rect 919 121 921 123
rect 889 108 891 110
rect 984 116 986 118
rect 903 108 905 110
rect 1024 116 1026 118
rect 994 109 996 111
rect 1064 121 1066 123
rect 1034 108 1036 110
rect 1129 116 1131 118
rect 1048 108 1050 110
rect 1169 121 1171 123
rect 1139 108 1141 110
rect 1153 108 1155 110
rect 36 43 38 45
rect 26 36 28 38
rect 76 44 78 46
rect 90 44 92 46
rect 66 36 68 38
rect 181 44 183 46
rect 195 44 197 46
rect 106 31 108 33
rect 171 36 173 38
rect 286 43 288 45
rect 211 31 213 33
rect 276 36 278 38
rect 326 44 328 46
rect 340 44 342 46
rect 316 36 318 38
rect 431 44 433 46
rect 445 44 447 46
rect 356 31 358 33
rect 421 36 423 38
rect 536 43 538 45
rect 461 31 463 33
rect 526 36 528 38
rect 576 44 578 46
rect 590 44 592 46
rect 566 36 568 38
rect 681 44 683 46
rect 695 44 697 46
rect 606 31 608 33
rect 671 36 673 38
rect 786 43 788 45
rect 711 31 713 33
rect 776 36 778 38
rect 826 44 828 46
rect 840 44 842 46
rect 816 36 818 38
rect 931 44 933 46
rect 945 44 947 46
rect 856 31 858 33
rect 921 36 923 38
rect 961 31 963 33
<< ndifct0 >>
rect 16 401 18 403
rect 56 401 58 403
rect 131 399 133 401
rect 143 402 145 404
rect 168 401 170 403
rect 157 394 159 396
rect 498 403 500 405
rect 538 403 540 405
rect 613 401 615 403
rect 625 404 627 406
rect 650 403 652 405
rect 639 396 641 398
rect 703 403 705 405
rect 743 403 745 405
rect 818 401 820 403
rect 830 404 832 406
rect 855 403 857 405
rect 844 396 846 398
rect 46 289 48 291
rect 56 289 58 291
rect 137 296 139 298
rect 126 289 128 291
rect 151 288 153 290
rect 163 291 165 293
rect 528 291 530 293
rect 538 291 540 293
rect 619 298 621 300
rect 608 291 610 293
rect 633 290 635 292
rect 645 293 647 295
rect 733 291 735 293
rect 743 291 745 293
rect 824 298 826 300
rect 813 291 815 293
rect 838 290 840 292
rect 850 293 852 295
rect 1024 285 1026 287
rect 1064 285 1066 287
rect 1139 283 1141 285
rect 1151 286 1153 288
rect 1176 285 1178 287
rect 1165 278 1167 280
rect 23 180 25 182
rect 14 167 16 169
rect 84 180 86 182
rect 73 173 75 175
rect 98 172 100 174
rect 33 167 35 169
rect 110 175 112 177
rect 189 180 191 182
rect 178 173 180 175
rect 203 172 205 174
rect 215 175 217 177
rect 273 180 275 182
rect 264 167 266 169
rect 334 180 336 182
rect 323 173 325 175
rect 348 172 350 174
rect 283 167 285 169
rect 360 175 362 177
rect 439 180 441 182
rect 428 173 430 175
rect 453 172 455 174
rect 465 175 467 177
rect 523 180 525 182
rect 514 167 516 169
rect 584 180 586 182
rect 573 173 575 175
rect 598 172 600 174
rect 533 167 535 169
rect 610 175 612 177
rect 689 180 691 182
rect 678 173 680 175
rect 703 172 705 174
rect 715 175 717 177
rect 773 180 775 182
rect 764 167 766 169
rect 834 180 836 182
rect 823 173 825 175
rect 848 172 850 174
rect 783 167 785 169
rect 860 175 862 177
rect 939 180 941 182
rect 928 173 930 175
rect 953 172 955 174
rect 965 175 967 177
rect 1054 173 1056 175
rect 1064 173 1066 175
rect 1145 180 1147 182
rect 1134 173 1136 175
rect 1159 172 1161 174
rect 1171 175 1173 177
rect 132 132 134 134
rect 157 133 159 135
rect 143 125 145 127
rect 169 130 171 132
rect 228 138 230 140
rect 247 138 249 140
rect 237 125 239 127
rect 287 132 289 134
rect 312 133 314 135
rect 298 125 300 127
rect 324 130 326 132
rect 392 132 394 134
rect 417 133 419 135
rect 403 125 405 127
rect 429 130 431 132
rect 478 138 480 140
rect 497 138 499 140
rect 487 125 489 127
rect 537 132 539 134
rect 562 133 564 135
rect 548 125 550 127
rect 574 130 576 132
rect 642 132 644 134
rect 667 133 669 135
rect 653 125 655 127
rect 679 130 681 132
rect 728 138 730 140
rect 747 138 749 140
rect 737 125 739 127
rect 787 132 789 134
rect 812 133 814 135
rect 798 125 800 127
rect 824 130 826 132
rect 892 132 894 134
rect 917 133 919 135
rect 903 125 905 127
rect 929 130 931 132
rect 978 138 980 140
rect 997 138 999 140
rect 987 125 989 127
rect 1037 132 1039 134
rect 1062 133 1064 135
rect 1048 125 1050 127
rect 1074 130 1076 132
rect 1142 132 1144 134
rect 1167 133 1169 135
rect 1153 125 1155 127
rect 1179 130 1181 132
rect 29 27 31 29
rect 20 14 22 16
rect 90 27 92 29
rect 79 20 81 22
rect 104 19 106 21
rect 39 14 41 16
rect 116 22 118 24
rect 195 27 197 29
rect 184 20 186 22
rect 209 19 211 21
rect 221 22 223 24
rect 279 27 281 29
rect 270 14 272 16
rect 340 27 342 29
rect 329 20 331 22
rect 354 19 356 21
rect 289 14 291 16
rect 366 22 368 24
rect 445 27 447 29
rect 434 20 436 22
rect 459 19 461 21
rect 471 22 473 24
rect 529 27 531 29
rect 520 14 522 16
rect 590 27 592 29
rect 579 20 581 22
rect 604 19 606 21
rect 539 14 541 16
rect 616 22 618 24
rect 695 27 697 29
rect 684 20 686 22
rect 709 19 711 21
rect 721 22 723 24
rect 779 27 781 29
rect 770 14 772 16
rect 840 27 842 29
rect 829 20 831 22
rect 854 19 856 21
rect 789 14 791 16
rect 866 22 868 24
rect 945 27 947 29
rect 934 20 936 22
rect 959 19 961 21
rect 971 22 973 24
<< ndifct1 >>
rect 35 411 37 413
rect 75 411 77 413
rect 103 411 105 413
rect 46 399 48 401
rect 86 399 88 401
rect 187 411 189 413
rect 121 401 123 403
rect 517 413 519 415
rect 557 413 559 415
rect 198 399 200 401
rect 585 413 587 415
rect 528 401 530 403
rect 568 401 570 403
rect 669 413 671 415
rect 603 403 605 405
rect 722 413 724 415
rect 762 413 764 415
rect 680 401 682 403
rect 790 413 792 415
rect 733 401 735 403
rect 773 401 775 403
rect 874 413 876 415
rect 808 403 810 405
rect 885 401 887 403
rect 16 291 18 293
rect 86 291 88 293
rect 96 291 98 293
rect 27 279 29 281
rect 75 279 77 281
rect 173 289 175 291
rect 107 279 109 281
rect 498 293 500 295
rect 568 293 570 295
rect 578 293 580 295
rect 191 279 193 281
rect 509 281 511 283
rect 557 281 559 283
rect 655 291 657 293
rect 589 281 591 283
rect 703 293 705 295
rect 773 293 775 295
rect 783 293 785 295
rect 673 281 675 283
rect 714 281 716 283
rect 762 281 764 283
rect 860 291 862 293
rect 794 281 796 283
rect 1043 295 1045 297
rect 1083 295 1085 297
rect 878 281 880 283
rect 1111 295 1113 297
rect 1054 283 1056 285
rect 1094 283 1096 285
rect 1195 295 1197 297
rect 1129 285 1131 287
rect 1206 283 1208 285
rect 3 180 5 182
rect 43 175 45 177
rect 120 173 122 175
rect 54 163 56 165
rect 148 175 150 177
rect 253 180 255 182
rect 138 163 140 165
rect 225 173 227 175
rect 159 163 161 165
rect 293 175 295 177
rect 243 163 245 165
rect 370 173 372 175
rect 304 163 306 165
rect 398 175 400 177
rect 503 180 505 182
rect 388 163 390 165
rect 475 173 477 175
rect 409 163 411 165
rect 543 175 545 177
rect 493 163 495 165
rect 620 173 622 175
rect 554 163 556 165
rect 648 175 650 177
rect 753 180 755 182
rect 638 163 640 165
rect 725 173 727 175
rect 659 163 661 165
rect 793 175 795 177
rect 743 163 745 165
rect 870 173 872 175
rect 804 163 806 165
rect 898 175 900 177
rect 888 163 890 165
rect 975 173 977 175
rect 909 163 911 165
rect 1024 175 1026 177
rect 1094 175 1096 177
rect 1104 175 1106 177
rect 993 163 995 165
rect 1035 163 1037 165
rect 1083 163 1085 165
rect 1181 173 1183 175
rect 1115 163 1117 165
rect 1199 163 1201 165
rect 113 142 115 144
rect 197 142 199 144
rect 102 130 104 132
rect 179 132 181 134
rect 268 142 270 144
rect 217 125 219 127
rect 352 142 354 144
rect 373 142 375 144
rect 257 130 259 132
rect 334 132 336 134
rect 457 142 459 144
rect 362 130 364 132
rect 439 132 441 134
rect 518 142 520 144
rect 467 125 469 127
rect 602 142 604 144
rect 623 142 625 144
rect 507 130 509 132
rect 584 132 586 134
rect 707 142 709 144
rect 612 130 614 132
rect 689 132 691 134
rect 768 142 770 144
rect 717 125 719 127
rect 852 142 854 144
rect 873 142 875 144
rect 757 130 759 132
rect 834 132 836 134
rect 957 142 959 144
rect 862 130 864 132
rect 939 132 941 134
rect 1018 142 1020 144
rect 967 125 969 127
rect 1102 142 1104 144
rect 1123 142 1125 144
rect 1007 130 1009 132
rect 1084 132 1086 134
rect 1207 142 1209 144
rect 1112 130 1114 132
rect 1189 132 1191 134
rect 9 27 11 29
rect 49 22 51 24
rect 126 20 128 22
rect 60 10 62 12
rect 154 22 156 24
rect 259 27 261 29
rect 144 10 146 12
rect 231 20 233 22
rect 165 10 167 12
rect 299 22 301 24
rect 249 10 251 12
rect 376 20 378 22
rect 310 10 312 12
rect 404 22 406 24
rect 509 27 511 29
rect 394 10 396 12
rect 481 20 483 22
rect 415 10 417 12
rect 549 22 551 24
rect 499 10 501 12
rect 626 20 628 22
rect 560 10 562 12
rect 654 22 656 24
rect 759 27 761 29
rect 644 10 646 12
rect 731 20 733 22
rect 665 10 667 12
rect 799 22 801 24
rect 749 10 751 12
rect 876 20 878 22
rect 810 10 812 12
rect 904 22 906 24
rect 894 10 896 12
rect 981 20 983 22
rect 915 10 917 12
rect 999 10 1001 12
<< ntiect1 >>
rect 45 351 47 353
rect 85 351 87 353
rect 123 351 125 353
rect 197 351 199 353
rect 527 353 529 355
rect 567 353 569 355
rect 605 353 607 355
rect 679 353 681 355
rect 732 353 734 355
rect 772 353 774 355
rect 810 353 812 355
rect 884 353 886 355
rect 17 339 19 341
rect 85 339 87 341
rect 97 339 99 341
rect 171 339 173 341
rect 499 341 501 343
rect 567 341 569 343
rect 579 341 581 343
rect 653 341 655 343
rect 704 341 706 343
rect 772 341 774 343
rect 784 341 786 343
rect 858 341 860 343
rect 1053 235 1055 237
rect 1093 235 1095 237
rect 1131 235 1133 237
rect 1205 235 1207 237
rect 4 223 6 225
rect 44 223 46 225
rect 118 223 120 225
rect 149 223 151 225
rect 223 223 225 225
rect 254 223 256 225
rect 294 223 296 225
rect 368 223 370 225
rect 399 223 401 225
rect 473 223 475 225
rect 504 223 506 225
rect 544 223 546 225
rect 618 223 620 225
rect 649 223 651 225
rect 723 223 725 225
rect 754 223 756 225
rect 794 223 796 225
rect 868 223 870 225
rect 899 223 901 225
rect 973 223 975 225
rect 1025 223 1027 225
rect 1093 223 1095 225
rect 1105 223 1107 225
rect 1179 223 1181 225
rect 103 82 105 84
rect 177 82 179 84
rect 218 82 220 84
rect 258 82 260 84
rect 332 82 334 84
rect 363 82 365 84
rect 437 82 439 84
rect 468 82 470 84
rect 508 82 510 84
rect 582 82 584 84
rect 613 82 615 84
rect 687 82 689 84
rect 718 82 720 84
rect 758 82 760 84
rect 832 82 834 84
rect 863 82 865 84
rect 937 82 939 84
rect 968 82 970 84
rect 1008 82 1010 84
rect 1082 82 1084 84
rect 1113 82 1115 84
rect 1187 82 1189 84
rect 10 70 12 72
rect 50 70 52 72
rect 124 70 126 72
rect 155 70 157 72
rect 229 70 231 72
rect 260 70 262 72
rect 300 70 302 72
rect 374 70 376 72
rect 405 70 407 72
rect 479 70 481 72
rect 510 70 512 72
rect 550 70 552 72
rect 624 70 626 72
rect 655 70 657 72
rect 729 70 731 72
rect 760 70 762 72
rect 800 70 802 72
rect 874 70 876 72
rect 905 70 907 72
rect 979 70 981 72
<< ptiect1 >>
rect 45 411 47 413
rect 85 411 87 413
rect 156 411 158 413
rect 197 411 199 413
rect 527 413 529 415
rect 567 413 569 415
rect 638 413 640 415
rect 679 413 681 415
rect 732 413 734 415
rect 772 413 774 415
rect 843 413 845 415
rect 884 413 886 415
rect 17 279 19 281
rect 85 279 87 281
rect 97 279 99 281
rect 138 279 140 281
rect 499 281 501 283
rect 567 281 569 283
rect 579 281 581 283
rect 620 281 622 283
rect 704 281 706 283
rect 772 281 774 283
rect 784 281 786 283
rect 825 281 827 283
rect 1053 295 1055 297
rect 1093 295 1095 297
rect 1164 295 1166 297
rect 1205 295 1207 297
rect 4 163 6 165
rect 44 163 46 165
rect 85 163 87 165
rect 149 163 151 165
rect 190 163 192 165
rect 254 163 256 165
rect 294 163 296 165
rect 335 163 337 165
rect 399 163 401 165
rect 440 163 442 165
rect 504 163 506 165
rect 544 163 546 165
rect 585 163 587 165
rect 649 163 651 165
rect 690 163 692 165
rect 754 163 756 165
rect 794 163 796 165
rect 835 163 837 165
rect 899 163 901 165
rect 940 163 942 165
rect 1025 163 1027 165
rect 1093 163 1095 165
rect 1105 163 1107 165
rect 1146 163 1148 165
rect 103 142 105 144
rect 144 142 146 144
rect 218 142 220 144
rect 258 142 260 144
rect 299 142 301 144
rect 363 142 365 144
rect 404 142 406 144
rect 468 142 470 144
rect 508 142 510 144
rect 549 142 551 144
rect 613 142 615 144
rect 654 142 656 144
rect 718 142 720 144
rect 758 142 760 144
rect 799 142 801 144
rect 863 142 865 144
rect 904 142 906 144
rect 968 142 970 144
rect 1008 142 1010 144
rect 1049 142 1051 144
rect 1113 142 1115 144
rect 1154 142 1156 144
rect 10 10 12 12
rect 50 10 52 12
rect 91 10 93 12
rect 155 10 157 12
rect 196 10 198 12
rect 260 10 262 12
rect 300 10 302 12
rect 341 10 343 12
rect 405 10 407 12
rect 446 10 448 12
rect 510 10 512 12
rect 550 10 552 12
rect 591 10 593 12
rect 655 10 657 12
rect 696 10 698 12
rect 760 10 762 12
rect 800 10 802 12
rect 841 10 843 12
rect 905 10 907 12
rect 946 10 948 12
<< pdifct0 >>
rect 16 361 18 363
rect 26 368 28 370
rect 26 361 28 363
rect 36 363 38 365
rect 56 361 58 363
rect 66 368 68 370
rect 66 361 68 363
rect 76 363 78 365
rect 103 360 105 362
rect 123 375 125 377
rect 123 368 125 370
rect 139 361 141 363
rect 139 354 141 356
rect 149 375 151 377
rect 168 361 170 363
rect 178 368 180 370
rect 178 361 180 363
rect 188 363 190 365
rect 498 363 500 365
rect 508 370 510 372
rect 508 363 510 365
rect 518 365 520 367
rect 538 363 540 365
rect 548 370 550 372
rect 548 363 550 365
rect 558 365 560 367
rect 585 362 587 364
rect 605 377 607 379
rect 605 370 607 372
rect 621 363 623 365
rect 621 356 623 358
rect 631 377 633 379
rect 650 363 652 365
rect 660 370 662 372
rect 660 363 662 365
rect 670 365 672 367
rect 703 363 705 365
rect 713 370 715 372
rect 713 363 715 365
rect 723 365 725 367
rect 743 363 745 365
rect 753 370 755 372
rect 753 363 755 365
rect 763 365 765 367
rect 790 362 792 364
rect 810 377 812 379
rect 810 370 812 372
rect 826 363 828 365
rect 826 356 828 358
rect 836 377 838 379
rect 855 363 857 365
rect 865 370 867 372
rect 865 363 867 365
rect 875 365 877 367
rect 26 327 28 329
rect 36 329 38 331
rect 36 322 38 324
rect 46 329 48 331
rect 56 329 58 331
rect 66 329 68 331
rect 66 322 68 324
rect 76 327 78 329
rect 106 327 108 329
rect 116 329 118 331
rect 116 322 118 324
rect 126 329 128 331
rect 145 315 147 317
rect 155 336 157 338
rect 155 329 157 331
rect 171 322 173 324
rect 171 315 173 317
rect 191 330 193 332
rect 508 329 510 331
rect 518 331 520 333
rect 518 324 520 326
rect 528 331 530 333
rect 538 331 540 333
rect 548 331 550 333
rect 548 324 550 326
rect 558 329 560 331
rect 588 329 590 331
rect 598 331 600 333
rect 598 324 600 326
rect 608 331 610 333
rect 627 317 629 319
rect 637 338 639 340
rect 637 331 639 333
rect 653 324 655 326
rect 653 317 655 319
rect 673 332 675 334
rect 713 329 715 331
rect 723 331 725 333
rect 723 324 725 326
rect 733 331 735 333
rect 743 331 745 333
rect 753 331 755 333
rect 753 324 755 326
rect 763 329 765 331
rect 793 329 795 331
rect 803 331 805 333
rect 803 324 805 326
rect 813 331 815 333
rect 832 317 834 319
rect 842 338 844 340
rect 842 331 844 333
rect 858 324 860 326
rect 858 317 860 319
rect 878 332 880 334
rect 1024 245 1026 247
rect 1034 252 1036 254
rect 1034 245 1036 247
rect 1044 247 1046 249
rect 1064 245 1066 247
rect 1074 252 1076 254
rect 1074 245 1076 247
rect 1084 247 1086 249
rect 1111 244 1113 246
rect 1131 259 1133 261
rect 1131 252 1133 254
rect 1147 245 1149 247
rect 1147 238 1149 240
rect 1157 259 1159 261
rect 1176 245 1178 247
rect 1186 252 1188 254
rect 1186 245 1188 247
rect 1196 247 1198 249
rect 14 220 16 222
rect 33 213 35 215
rect 53 211 55 213
rect 63 213 65 215
rect 63 206 65 208
rect 73 213 75 215
rect 92 199 94 201
rect 102 220 104 222
rect 102 213 104 215
rect 118 206 120 208
rect 118 199 120 201
rect 138 214 140 216
rect 158 211 160 213
rect 168 213 170 215
rect 168 206 170 208
rect 178 213 180 215
rect 197 199 199 201
rect 207 220 209 222
rect 207 213 209 215
rect 223 206 225 208
rect 223 199 225 201
rect 264 220 266 222
rect 243 214 245 216
rect 283 213 285 215
rect 303 211 305 213
rect 313 213 315 215
rect 313 206 315 208
rect 323 213 325 215
rect 342 199 344 201
rect 352 220 354 222
rect 352 213 354 215
rect 368 206 370 208
rect 368 199 370 201
rect 388 214 390 216
rect 408 211 410 213
rect 418 213 420 215
rect 418 206 420 208
rect 428 213 430 215
rect 447 199 449 201
rect 457 220 459 222
rect 457 213 459 215
rect 473 206 475 208
rect 473 199 475 201
rect 514 220 516 222
rect 493 214 495 216
rect 533 213 535 215
rect 553 211 555 213
rect 563 213 565 215
rect 563 206 565 208
rect 573 213 575 215
rect 592 199 594 201
rect 602 220 604 222
rect 602 213 604 215
rect 618 206 620 208
rect 618 199 620 201
rect 638 214 640 216
rect 658 211 660 213
rect 668 213 670 215
rect 668 206 670 208
rect 678 213 680 215
rect 697 199 699 201
rect 707 220 709 222
rect 707 213 709 215
rect 723 206 725 208
rect 723 199 725 201
rect 764 220 766 222
rect 743 214 745 216
rect 783 213 785 215
rect 803 211 805 213
rect 813 213 815 215
rect 813 206 815 208
rect 823 213 825 215
rect 842 199 844 201
rect 852 220 854 222
rect 852 213 854 215
rect 868 206 870 208
rect 868 199 870 201
rect 888 214 890 216
rect 908 211 910 213
rect 918 213 920 215
rect 918 206 920 208
rect 928 213 930 215
rect 947 199 949 201
rect 957 220 959 222
rect 957 213 959 215
rect 973 206 975 208
rect 973 199 975 201
rect 993 214 995 216
rect 1034 211 1036 213
rect 1044 213 1046 215
rect 1044 206 1046 208
rect 1054 213 1056 215
rect 1064 213 1066 215
rect 1074 213 1076 215
rect 1074 206 1076 208
rect 1084 211 1086 213
rect 1114 211 1116 213
rect 1124 213 1126 215
rect 1124 206 1126 208
rect 1134 213 1136 215
rect 1153 199 1155 201
rect 1163 220 1165 222
rect 1163 213 1165 215
rect 1179 206 1181 208
rect 1179 199 1181 201
rect 1199 214 1201 216
rect 151 106 153 108
rect 112 94 114 96
rect 122 99 124 101
rect 122 92 124 94
rect 132 92 134 94
rect 161 92 163 94
rect 177 106 179 108
rect 177 99 179 101
rect 161 85 163 87
rect 197 91 199 93
rect 228 85 230 87
rect 247 92 249 94
rect 306 106 308 108
rect 267 94 269 96
rect 277 99 279 101
rect 277 92 279 94
rect 287 92 289 94
rect 316 92 318 94
rect 332 106 334 108
rect 332 99 334 101
rect 316 85 318 87
rect 352 91 354 93
rect 411 106 413 108
rect 372 94 374 96
rect 382 99 384 101
rect 382 92 384 94
rect 392 92 394 94
rect 421 92 423 94
rect 437 106 439 108
rect 437 99 439 101
rect 421 85 423 87
rect 457 91 459 93
rect 478 85 480 87
rect 497 92 499 94
rect 556 106 558 108
rect 517 94 519 96
rect 527 99 529 101
rect 527 92 529 94
rect 537 92 539 94
rect 566 92 568 94
rect 582 106 584 108
rect 582 99 584 101
rect 566 85 568 87
rect 602 91 604 93
rect 661 106 663 108
rect 622 94 624 96
rect 632 99 634 101
rect 632 92 634 94
rect 642 92 644 94
rect 671 92 673 94
rect 687 106 689 108
rect 687 99 689 101
rect 671 85 673 87
rect 707 91 709 93
rect 728 85 730 87
rect 747 92 749 94
rect 806 106 808 108
rect 767 94 769 96
rect 777 99 779 101
rect 777 92 779 94
rect 787 92 789 94
rect 816 92 818 94
rect 832 106 834 108
rect 832 99 834 101
rect 816 85 818 87
rect 852 91 854 93
rect 911 106 913 108
rect 872 94 874 96
rect 882 99 884 101
rect 882 92 884 94
rect 892 92 894 94
rect 921 92 923 94
rect 937 106 939 108
rect 937 99 939 101
rect 921 85 923 87
rect 957 91 959 93
rect 978 85 980 87
rect 997 92 999 94
rect 1056 106 1058 108
rect 1017 94 1019 96
rect 1027 99 1029 101
rect 1027 92 1029 94
rect 1037 92 1039 94
rect 1066 92 1068 94
rect 1082 106 1084 108
rect 1082 99 1084 101
rect 1066 85 1068 87
rect 1102 91 1104 93
rect 1161 106 1163 108
rect 1122 94 1124 96
rect 1132 99 1134 101
rect 1132 92 1134 94
rect 1142 92 1144 94
rect 1171 92 1173 94
rect 1187 106 1189 108
rect 1187 99 1189 101
rect 1171 85 1173 87
rect 1207 91 1209 93
rect 20 67 22 69
rect 39 60 41 62
rect 59 58 61 60
rect 69 60 71 62
rect 69 53 71 55
rect 79 60 81 62
rect 98 46 100 48
rect 108 67 110 69
rect 108 60 110 62
rect 124 53 126 55
rect 124 46 126 48
rect 144 61 146 63
rect 164 58 166 60
rect 174 60 176 62
rect 174 53 176 55
rect 184 60 186 62
rect 203 46 205 48
rect 213 67 215 69
rect 213 60 215 62
rect 229 53 231 55
rect 229 46 231 48
rect 270 67 272 69
rect 249 61 251 63
rect 289 60 291 62
rect 309 58 311 60
rect 319 60 321 62
rect 319 53 321 55
rect 329 60 331 62
rect 348 46 350 48
rect 358 67 360 69
rect 358 60 360 62
rect 374 53 376 55
rect 374 46 376 48
rect 394 61 396 63
rect 414 58 416 60
rect 424 60 426 62
rect 424 53 426 55
rect 434 60 436 62
rect 453 46 455 48
rect 463 67 465 69
rect 463 60 465 62
rect 479 53 481 55
rect 479 46 481 48
rect 520 67 522 69
rect 499 61 501 63
rect 539 60 541 62
rect 559 58 561 60
rect 569 60 571 62
rect 569 53 571 55
rect 579 60 581 62
rect 598 46 600 48
rect 608 67 610 69
rect 608 60 610 62
rect 624 53 626 55
rect 624 46 626 48
rect 644 61 646 63
rect 664 58 666 60
rect 674 60 676 62
rect 674 53 676 55
rect 684 60 686 62
rect 703 46 705 48
rect 713 67 715 69
rect 713 60 715 62
rect 729 53 731 55
rect 729 46 731 48
rect 770 67 772 69
rect 749 61 751 63
rect 789 60 791 62
rect 809 58 811 60
rect 819 60 821 62
rect 819 53 821 55
rect 829 60 831 62
rect 848 46 850 48
rect 858 67 860 69
rect 858 60 860 62
rect 874 53 876 55
rect 874 46 876 48
rect 894 61 896 63
rect 914 58 916 60
rect 924 60 926 62
rect 924 53 926 55
rect 934 60 936 62
rect 953 46 955 48
rect 963 67 965 69
rect 963 60 965 62
rect 979 53 981 55
rect 979 46 981 48
rect 999 61 1001 63
<< pdifct1 >>
rect 46 375 48 377
rect 46 368 48 370
rect 86 375 88 377
rect 86 368 88 370
rect 113 368 115 370
rect 198 375 200 377
rect 198 368 200 370
rect 528 377 530 379
rect 528 370 530 372
rect 568 377 570 379
rect 568 370 570 372
rect 595 370 597 372
rect 680 377 682 379
rect 680 370 682 372
rect 733 377 735 379
rect 733 370 735 372
rect 773 377 775 379
rect 773 370 775 372
rect 800 370 802 372
rect 885 377 887 379
rect 885 370 887 372
rect 16 322 18 324
rect 16 315 18 317
rect 86 322 88 324
rect 86 315 88 317
rect 96 322 98 324
rect 96 315 98 317
rect 181 322 183 324
rect 498 324 500 326
rect 498 317 500 319
rect 568 324 570 326
rect 568 317 570 319
rect 578 324 580 326
rect 578 317 580 319
rect 663 324 665 326
rect 703 324 705 326
rect 703 317 705 319
rect 773 324 775 326
rect 773 317 775 319
rect 783 324 785 326
rect 783 317 785 319
rect 868 324 870 326
rect 1054 259 1056 261
rect 1054 252 1056 254
rect 1094 259 1096 261
rect 1094 252 1096 254
rect 1121 252 1123 254
rect 1206 259 1208 261
rect 1206 252 1208 254
rect 3 210 5 212
rect 3 203 5 205
rect 43 206 45 208
rect 43 199 45 201
rect 128 206 130 208
rect 148 206 150 208
rect 148 199 150 201
rect 233 206 235 208
rect 253 210 255 212
rect 253 203 255 205
rect 293 206 295 208
rect 293 199 295 201
rect 378 206 380 208
rect 398 206 400 208
rect 398 199 400 201
rect 483 206 485 208
rect 503 210 505 212
rect 503 203 505 205
rect 543 206 545 208
rect 543 199 545 201
rect 628 206 630 208
rect 648 206 650 208
rect 648 199 650 201
rect 733 206 735 208
rect 753 210 755 212
rect 753 203 755 205
rect 793 206 795 208
rect 793 199 795 201
rect 878 206 880 208
rect 898 206 900 208
rect 898 199 900 201
rect 983 206 985 208
rect 1024 206 1026 208
rect 1024 199 1026 201
rect 1094 206 1096 208
rect 1094 199 1096 201
rect 1104 206 1106 208
rect 1104 199 1106 201
rect 1189 206 1191 208
rect 102 106 104 108
rect 102 99 104 101
rect 187 99 189 101
rect 217 102 219 104
rect 217 95 219 97
rect 257 106 259 108
rect 257 99 259 101
rect 342 99 344 101
rect 362 106 364 108
rect 362 99 364 101
rect 447 99 449 101
rect 467 102 469 104
rect 467 95 469 97
rect 507 106 509 108
rect 507 99 509 101
rect 592 99 594 101
rect 612 106 614 108
rect 612 99 614 101
rect 697 99 699 101
rect 717 102 719 104
rect 717 95 719 97
rect 757 106 759 108
rect 757 99 759 101
rect 842 99 844 101
rect 862 106 864 108
rect 862 99 864 101
rect 947 99 949 101
rect 967 102 969 104
rect 967 95 969 97
rect 1007 106 1009 108
rect 1007 99 1009 101
rect 1092 99 1094 101
rect 1112 106 1114 108
rect 1112 99 1114 101
rect 1197 99 1199 101
rect 9 57 11 59
rect 9 50 11 52
rect 49 53 51 55
rect 49 46 51 48
rect 134 53 136 55
rect 154 53 156 55
rect 154 46 156 48
rect 239 53 241 55
rect 259 57 261 59
rect 259 50 261 52
rect 299 53 301 55
rect 299 46 301 48
rect 384 53 386 55
rect 404 53 406 55
rect 404 46 406 48
rect 489 53 491 55
rect 509 57 511 59
rect 509 50 511 52
rect 549 53 551 55
rect 549 46 551 48
rect 634 53 636 55
rect 654 53 656 55
rect 654 46 656 48
rect 739 53 741 55
rect 759 57 761 59
rect 759 50 761 52
rect 799 53 801 55
rect 799 46 801 48
rect 884 53 886 55
rect 904 53 906 55
rect 904 46 906 48
rect 989 53 991 55
<< alu0 >>
rect 14 403 34 404
rect 14 401 16 403
rect 18 401 34 403
rect 14 400 34 401
rect 30 396 34 400
rect 54 403 74 404
rect 54 401 56 403
rect 58 401 74 403
rect 54 400 74 401
rect 45 397 46 399
rect 30 392 42 396
rect 38 387 42 392
rect 38 385 39 387
rect 41 385 42 387
rect 38 373 42 385
rect 70 396 74 400
rect 141 404 147 410
rect 496 405 516 406
rect 85 397 86 399
rect 70 392 82 396
rect 78 387 82 392
rect 78 385 79 387
rect 81 385 82 387
rect 25 370 42 373
rect 25 368 26 370
rect 28 369 42 370
rect 28 368 29 369
rect 14 363 20 364
rect 14 361 16 363
rect 18 361 20 363
rect 14 354 20 361
rect 25 363 29 368
rect 78 373 82 385
rect 65 370 82 373
rect 65 368 66 370
rect 68 369 82 370
rect 68 368 69 369
rect 25 361 26 363
rect 28 361 29 363
rect 25 359 29 361
rect 34 365 40 366
rect 34 363 36 365
rect 38 363 40 365
rect 34 354 40 363
rect 54 363 60 364
rect 54 361 56 363
rect 58 361 60 363
rect 54 354 60 361
rect 65 363 69 368
rect 130 401 134 403
rect 141 402 143 404
rect 145 402 147 404
rect 141 401 147 402
rect 166 403 186 404
rect 166 401 168 403
rect 170 401 186 403
rect 130 399 131 401
rect 133 399 134 401
rect 166 400 186 401
rect 130 396 134 399
rect 110 392 134 396
rect 110 388 114 392
rect 156 396 160 398
rect 156 394 157 396
rect 159 394 160 396
rect 109 386 114 388
rect 109 384 110 386
rect 112 384 114 386
rect 118 387 134 388
rect 118 385 120 387
rect 122 385 134 387
rect 118 384 134 385
rect 109 382 114 384
rect 110 380 114 382
rect 110 377 126 380
rect 110 376 123 377
rect 122 375 123 376
rect 125 375 126 377
rect 122 370 126 375
rect 122 368 123 370
rect 125 368 126 370
rect 122 366 126 368
rect 130 378 134 384
rect 156 388 160 394
rect 149 384 160 388
rect 182 396 186 400
rect 496 403 498 405
rect 500 403 516 405
rect 496 402 516 403
rect 197 397 198 399
rect 182 392 194 396
rect 190 387 194 392
rect 190 385 191 387
rect 193 385 194 387
rect 149 378 153 384
rect 130 377 153 378
rect 130 375 149 377
rect 151 375 153 377
rect 130 374 153 375
rect 65 361 66 363
rect 68 361 69 363
rect 65 359 69 361
rect 74 365 80 366
rect 74 363 76 365
rect 78 363 80 365
rect 130 363 134 374
rect 190 373 194 385
rect 512 398 516 402
rect 536 405 556 406
rect 536 403 538 405
rect 540 403 556 405
rect 536 402 556 403
rect 527 399 528 401
rect 512 394 524 398
rect 520 389 524 394
rect 520 387 521 389
rect 523 387 524 389
rect 177 370 194 373
rect 177 368 178 370
rect 180 369 194 370
rect 180 368 181 369
rect 74 354 80 363
rect 101 362 134 363
rect 101 360 103 362
rect 105 360 134 362
rect 101 359 134 360
rect 138 363 142 365
rect 138 361 139 363
rect 141 361 142 363
rect 138 356 142 361
rect 166 363 172 364
rect 166 361 168 363
rect 170 361 172 363
rect 138 354 139 356
rect 141 354 142 356
rect 166 354 172 361
rect 177 363 181 368
rect 520 375 524 387
rect 552 398 556 402
rect 623 406 629 412
rect 567 399 568 401
rect 552 394 564 398
rect 560 389 564 394
rect 560 387 561 389
rect 563 387 564 389
rect 507 372 524 375
rect 507 370 508 372
rect 510 371 524 372
rect 510 370 511 371
rect 177 361 178 363
rect 180 361 181 363
rect 177 359 181 361
rect 186 365 192 366
rect 186 363 188 365
rect 190 363 192 365
rect 186 354 192 363
rect 496 365 502 366
rect 496 363 498 365
rect 500 363 502 365
rect 496 356 502 363
rect 507 365 511 370
rect 560 375 564 387
rect 547 372 564 375
rect 547 370 548 372
rect 550 371 564 372
rect 550 370 551 371
rect 507 363 508 365
rect 510 363 511 365
rect 507 361 511 363
rect 516 367 522 368
rect 516 365 518 367
rect 520 365 522 367
rect 516 356 522 365
rect 536 365 542 366
rect 536 363 538 365
rect 540 363 542 365
rect 536 356 542 363
rect 547 365 551 370
rect 612 403 616 405
rect 623 404 625 406
rect 627 404 629 406
rect 623 403 629 404
rect 648 405 668 406
rect 648 403 650 405
rect 652 403 668 405
rect 612 401 613 403
rect 615 401 616 403
rect 648 402 668 403
rect 612 398 616 401
rect 592 394 616 398
rect 592 390 596 394
rect 638 398 642 400
rect 638 396 639 398
rect 641 396 642 398
rect 591 388 596 390
rect 591 386 592 388
rect 594 386 596 388
rect 600 389 616 390
rect 600 387 602 389
rect 604 387 616 389
rect 600 386 616 387
rect 591 384 596 386
rect 592 382 596 384
rect 592 379 608 382
rect 592 378 605 379
rect 604 377 605 378
rect 607 377 608 379
rect 604 372 608 377
rect 604 370 605 372
rect 607 370 608 372
rect 604 368 608 370
rect 612 380 616 386
rect 638 390 642 396
rect 631 386 642 390
rect 664 398 668 402
rect 701 405 721 406
rect 701 403 703 405
rect 705 403 721 405
rect 701 402 721 403
rect 679 399 680 401
rect 664 394 676 398
rect 672 389 676 394
rect 672 387 673 389
rect 675 387 676 389
rect 631 380 635 386
rect 612 379 635 380
rect 612 377 631 379
rect 633 377 635 379
rect 612 376 635 377
rect 547 363 548 365
rect 550 363 551 365
rect 547 361 551 363
rect 556 367 562 368
rect 556 365 558 367
rect 560 365 562 367
rect 612 365 616 376
rect 672 375 676 387
rect 717 398 721 402
rect 741 405 761 406
rect 741 403 743 405
rect 745 403 761 405
rect 741 402 761 403
rect 732 399 733 401
rect 717 394 729 398
rect 725 389 729 394
rect 725 387 726 389
rect 728 387 729 389
rect 659 372 676 375
rect 659 370 660 372
rect 662 371 676 372
rect 662 370 663 371
rect 556 356 562 365
rect 583 364 616 365
rect 583 362 585 364
rect 587 362 616 364
rect 583 361 616 362
rect 620 365 624 367
rect 620 363 621 365
rect 623 363 624 365
rect 620 358 624 363
rect 648 365 654 366
rect 648 363 650 365
rect 652 363 654 365
rect 620 356 621 358
rect 623 356 624 358
rect 648 356 654 363
rect 659 365 663 370
rect 725 375 729 387
rect 757 398 761 402
rect 828 406 834 412
rect 772 399 773 401
rect 757 394 769 398
rect 765 389 769 394
rect 765 387 766 389
rect 768 387 769 389
rect 712 372 729 375
rect 712 370 713 372
rect 715 371 729 372
rect 715 370 716 371
rect 659 363 660 365
rect 662 363 663 365
rect 659 361 663 363
rect 668 367 674 368
rect 668 365 670 367
rect 672 365 674 367
rect 668 356 674 365
rect 701 365 707 366
rect 701 363 703 365
rect 705 363 707 365
rect 701 356 707 363
rect 712 365 716 370
rect 765 375 769 387
rect 752 372 769 375
rect 752 370 753 372
rect 755 371 769 372
rect 755 370 756 371
rect 712 363 713 365
rect 715 363 716 365
rect 712 361 716 363
rect 721 367 727 368
rect 721 365 723 367
rect 725 365 727 367
rect 721 356 727 365
rect 741 365 747 366
rect 741 363 743 365
rect 745 363 747 365
rect 741 356 747 363
rect 752 365 756 370
rect 817 403 821 405
rect 828 404 830 406
rect 832 404 834 406
rect 828 403 834 404
rect 853 405 873 406
rect 853 403 855 405
rect 857 403 873 405
rect 817 401 818 403
rect 820 401 821 403
rect 853 402 873 403
rect 817 398 821 401
rect 797 394 821 398
rect 797 390 801 394
rect 843 398 847 400
rect 843 396 844 398
rect 846 396 847 398
rect 796 388 801 390
rect 796 386 797 388
rect 799 386 801 388
rect 805 389 821 390
rect 805 387 807 389
rect 809 387 821 389
rect 805 386 821 387
rect 796 384 801 386
rect 797 382 801 384
rect 797 379 813 382
rect 797 378 810 379
rect 809 377 810 378
rect 812 377 813 379
rect 809 372 813 377
rect 809 370 810 372
rect 812 370 813 372
rect 809 368 813 370
rect 817 380 821 386
rect 843 390 847 396
rect 836 386 847 390
rect 869 398 873 402
rect 884 399 885 401
rect 869 394 881 398
rect 877 389 881 394
rect 877 387 878 389
rect 880 387 881 389
rect 836 380 840 386
rect 817 379 840 380
rect 817 377 836 379
rect 838 377 840 379
rect 817 376 840 377
rect 752 363 753 365
rect 755 363 756 365
rect 752 361 756 363
rect 761 367 767 368
rect 761 365 763 367
rect 765 365 767 367
rect 817 365 821 376
rect 877 375 881 387
rect 864 372 881 375
rect 864 370 865 372
rect 867 371 881 372
rect 867 370 868 371
rect 761 356 767 365
rect 788 364 821 365
rect 788 362 790 364
rect 792 362 821 364
rect 788 361 821 362
rect 825 365 829 367
rect 825 363 826 365
rect 828 363 829 365
rect 825 358 829 363
rect 853 365 859 366
rect 853 363 855 365
rect 857 363 859 365
rect 825 356 826 358
rect 828 356 829 358
rect 853 356 859 363
rect 864 365 868 370
rect 864 363 865 365
rect 867 363 868 365
rect 864 361 868 363
rect 873 367 879 368
rect 873 365 875 367
rect 877 365 879 367
rect 873 356 879 365
rect 24 329 30 338
rect 24 327 26 329
rect 28 327 30 329
rect 24 326 30 327
rect 35 331 39 333
rect 35 329 36 331
rect 38 329 39 331
rect 35 324 39 329
rect 44 331 50 338
rect 44 329 46 331
rect 48 329 50 331
rect 44 328 50 329
rect 54 331 60 338
rect 54 329 56 331
rect 58 329 60 331
rect 54 328 60 329
rect 65 331 69 333
rect 65 329 66 331
rect 68 329 69 331
rect 35 323 36 324
rect 22 322 36 323
rect 38 322 39 324
rect 22 319 39 322
rect 22 307 26 319
rect 65 324 69 329
rect 74 329 80 338
rect 74 327 76 329
rect 78 327 80 329
rect 74 326 80 327
rect 104 329 110 338
rect 104 327 106 329
rect 108 327 110 329
rect 104 326 110 327
rect 115 331 119 333
rect 115 329 116 331
rect 118 329 119 331
rect 65 322 66 324
rect 68 323 69 324
rect 68 322 82 323
rect 65 319 82 322
rect 22 305 23 307
rect 25 305 26 307
rect 22 300 26 305
rect 22 296 34 300
rect 18 293 19 295
rect 30 292 34 296
rect 78 307 82 319
rect 78 305 79 307
rect 81 305 82 307
rect 78 300 82 305
rect 70 296 82 300
rect 70 292 74 296
rect 85 293 86 295
rect 30 291 50 292
rect 30 289 46 291
rect 48 289 50 291
rect 30 288 50 289
rect 54 291 74 292
rect 54 289 56 291
rect 58 289 74 291
rect 54 288 74 289
rect 115 324 119 329
rect 124 331 130 338
rect 154 336 155 338
rect 157 336 158 338
rect 124 329 126 331
rect 128 329 130 331
rect 124 328 130 329
rect 154 331 158 336
rect 154 329 155 331
rect 157 329 158 331
rect 154 327 158 329
rect 162 332 195 333
rect 162 330 191 332
rect 193 330 195 332
rect 162 329 195 330
rect 506 331 512 340
rect 506 329 508 331
rect 510 329 512 331
rect 115 323 116 324
rect 102 322 116 323
rect 118 322 119 324
rect 102 319 119 322
rect 102 307 106 319
rect 162 318 166 329
rect 506 328 512 329
rect 517 333 521 335
rect 517 331 518 333
rect 520 331 521 333
rect 143 317 166 318
rect 143 315 145 317
rect 147 315 166 317
rect 143 314 166 315
rect 143 308 147 314
rect 102 305 103 307
rect 105 305 106 307
rect 102 300 106 305
rect 102 296 114 300
rect 98 293 99 295
rect 110 292 114 296
rect 136 304 147 308
rect 136 298 140 304
rect 162 308 166 314
rect 170 324 174 326
rect 170 322 171 324
rect 173 322 174 324
rect 170 317 174 322
rect 170 315 171 317
rect 173 316 174 317
rect 173 315 186 316
rect 170 312 186 315
rect 182 310 186 312
rect 182 308 187 310
rect 162 307 178 308
rect 162 305 174 307
rect 176 305 178 307
rect 162 304 178 305
rect 182 306 184 308
rect 186 306 187 308
rect 182 304 187 306
rect 136 296 137 298
rect 139 296 140 298
rect 136 294 140 296
rect 182 300 186 304
rect 162 296 186 300
rect 162 293 166 296
rect 110 291 130 292
rect 162 291 163 293
rect 165 291 166 293
rect 110 289 126 291
rect 128 289 130 291
rect 110 288 130 289
rect 149 290 155 291
rect 149 288 151 290
rect 153 288 155 290
rect 162 289 166 291
rect 517 326 521 331
rect 526 333 532 340
rect 526 331 528 333
rect 530 331 532 333
rect 526 330 532 331
rect 536 333 542 340
rect 536 331 538 333
rect 540 331 542 333
rect 536 330 542 331
rect 547 333 551 335
rect 547 331 548 333
rect 550 331 551 333
rect 517 325 518 326
rect 504 324 518 325
rect 520 324 521 326
rect 504 321 521 324
rect 504 309 508 321
rect 547 326 551 331
rect 556 331 562 340
rect 556 329 558 331
rect 560 329 562 331
rect 556 328 562 329
rect 586 331 592 340
rect 586 329 588 331
rect 590 329 592 331
rect 586 328 592 329
rect 597 333 601 335
rect 597 331 598 333
rect 600 331 601 333
rect 547 324 548 326
rect 550 325 551 326
rect 550 324 564 325
rect 547 321 564 324
rect 504 307 505 309
rect 507 307 508 309
rect 504 302 508 307
rect 504 298 516 302
rect 500 295 501 297
rect 512 294 516 298
rect 560 309 564 321
rect 560 307 561 309
rect 563 307 564 309
rect 560 302 564 307
rect 552 298 564 302
rect 552 294 556 298
rect 567 295 568 297
rect 512 293 532 294
rect 512 291 528 293
rect 530 291 532 293
rect 512 290 532 291
rect 536 293 556 294
rect 536 291 538 293
rect 540 291 556 293
rect 536 290 556 291
rect 597 326 601 331
rect 606 333 612 340
rect 636 338 637 340
rect 639 338 640 340
rect 606 331 608 333
rect 610 331 612 333
rect 606 330 612 331
rect 636 333 640 338
rect 636 331 637 333
rect 639 331 640 333
rect 636 329 640 331
rect 644 334 677 335
rect 644 332 673 334
rect 675 332 677 334
rect 644 331 677 332
rect 711 331 717 340
rect 597 325 598 326
rect 584 324 598 325
rect 600 324 601 326
rect 584 321 601 324
rect 584 309 588 321
rect 644 320 648 331
rect 711 329 713 331
rect 715 329 717 331
rect 711 328 717 329
rect 722 333 726 335
rect 722 331 723 333
rect 725 331 726 333
rect 625 319 648 320
rect 625 317 627 319
rect 629 317 648 319
rect 625 316 648 317
rect 625 310 629 316
rect 584 307 585 309
rect 587 307 588 309
rect 584 302 588 307
rect 584 298 596 302
rect 580 295 581 297
rect 592 294 596 298
rect 618 306 629 310
rect 618 300 622 306
rect 644 310 648 316
rect 652 326 656 328
rect 652 324 653 326
rect 655 324 656 326
rect 652 319 656 324
rect 652 317 653 319
rect 655 318 656 319
rect 655 317 668 318
rect 652 314 668 317
rect 664 312 668 314
rect 664 310 669 312
rect 644 309 660 310
rect 644 307 656 309
rect 658 307 660 309
rect 644 306 660 307
rect 664 308 666 310
rect 668 308 669 310
rect 664 306 669 308
rect 618 298 619 300
rect 621 298 622 300
rect 618 296 622 298
rect 664 302 668 306
rect 644 298 668 302
rect 644 295 648 298
rect 592 293 612 294
rect 644 293 645 295
rect 647 293 648 295
rect 592 291 608 293
rect 610 291 612 293
rect 592 290 612 291
rect 631 292 637 293
rect 631 290 633 292
rect 635 290 637 292
rect 644 291 648 293
rect 722 326 726 331
rect 731 333 737 340
rect 731 331 733 333
rect 735 331 737 333
rect 731 330 737 331
rect 741 333 747 340
rect 741 331 743 333
rect 745 331 747 333
rect 741 330 747 331
rect 752 333 756 335
rect 752 331 753 333
rect 755 331 756 333
rect 722 325 723 326
rect 709 324 723 325
rect 725 324 726 326
rect 709 321 726 324
rect 709 309 713 321
rect 752 326 756 331
rect 761 331 767 340
rect 761 329 763 331
rect 765 329 767 331
rect 761 328 767 329
rect 791 331 797 340
rect 791 329 793 331
rect 795 329 797 331
rect 791 328 797 329
rect 802 333 806 335
rect 802 331 803 333
rect 805 331 806 333
rect 752 324 753 326
rect 755 325 756 326
rect 755 324 769 325
rect 752 321 769 324
rect 709 307 710 309
rect 712 307 713 309
rect 709 302 713 307
rect 709 298 721 302
rect 705 295 706 297
rect 149 282 155 288
rect 631 284 637 290
rect 717 294 721 298
rect 765 309 769 321
rect 765 307 766 309
rect 768 307 769 309
rect 765 302 769 307
rect 757 298 769 302
rect 757 294 761 298
rect 772 295 773 297
rect 717 293 737 294
rect 717 291 733 293
rect 735 291 737 293
rect 717 290 737 291
rect 741 293 761 294
rect 741 291 743 293
rect 745 291 761 293
rect 741 290 761 291
rect 802 326 806 331
rect 811 333 817 340
rect 841 338 842 340
rect 844 338 845 340
rect 811 331 813 333
rect 815 331 817 333
rect 811 330 817 331
rect 841 333 845 338
rect 841 331 842 333
rect 844 331 845 333
rect 841 329 845 331
rect 849 334 882 335
rect 849 332 878 334
rect 880 332 882 334
rect 849 331 882 332
rect 802 325 803 326
rect 789 324 803 325
rect 805 324 806 326
rect 789 321 806 324
rect 789 309 793 321
rect 849 320 853 331
rect 830 319 853 320
rect 830 317 832 319
rect 834 317 853 319
rect 830 316 853 317
rect 830 310 834 316
rect 789 307 790 309
rect 792 307 793 309
rect 789 302 793 307
rect 789 298 801 302
rect 785 295 786 297
rect 797 294 801 298
rect 823 306 834 310
rect 823 300 827 306
rect 849 310 853 316
rect 857 326 861 328
rect 857 324 858 326
rect 860 324 861 326
rect 857 319 861 324
rect 857 317 858 319
rect 860 318 861 319
rect 860 317 873 318
rect 857 314 873 317
rect 869 312 873 314
rect 869 310 874 312
rect 849 309 865 310
rect 849 307 861 309
rect 863 307 865 309
rect 849 306 865 307
rect 869 308 871 310
rect 873 308 874 310
rect 869 306 874 308
rect 823 298 824 300
rect 826 298 827 300
rect 823 296 827 298
rect 869 302 873 306
rect 849 298 873 302
rect 849 295 853 298
rect 797 293 817 294
rect 849 293 850 295
rect 852 293 853 295
rect 797 291 813 293
rect 815 291 817 293
rect 797 290 817 291
rect 836 292 842 293
rect 836 290 838 292
rect 840 290 842 292
rect 849 291 853 293
rect 836 284 842 290
rect 1022 287 1042 288
rect 1022 285 1024 287
rect 1026 285 1042 287
rect 1022 284 1042 285
rect 1038 280 1042 284
rect 1062 287 1082 288
rect 1062 285 1064 287
rect 1066 285 1082 287
rect 1062 284 1082 285
rect 1053 281 1054 283
rect 1038 276 1050 280
rect 1046 271 1050 276
rect 1046 269 1047 271
rect 1049 269 1050 271
rect 1046 257 1050 269
rect 1078 280 1082 284
rect 1149 288 1155 294
rect 1093 281 1094 283
rect 1078 276 1090 280
rect 1086 271 1090 276
rect 1086 269 1087 271
rect 1089 269 1090 271
rect 1033 254 1050 257
rect 1033 252 1034 254
rect 1036 253 1050 254
rect 1036 252 1037 253
rect 1022 247 1028 248
rect 1022 245 1024 247
rect 1026 245 1028 247
rect 1022 238 1028 245
rect 1033 247 1037 252
rect 1086 257 1090 269
rect 1073 254 1090 257
rect 1073 252 1074 254
rect 1076 253 1090 254
rect 1076 252 1077 253
rect 1033 245 1034 247
rect 1036 245 1037 247
rect 1033 243 1037 245
rect 1042 249 1048 250
rect 1042 247 1044 249
rect 1046 247 1048 249
rect 1042 238 1048 247
rect 1062 247 1068 248
rect 1062 245 1064 247
rect 1066 245 1068 247
rect 1062 238 1068 245
rect 1073 247 1077 252
rect 1138 285 1142 287
rect 1149 286 1151 288
rect 1153 286 1155 288
rect 1149 285 1155 286
rect 1174 287 1194 288
rect 1174 285 1176 287
rect 1178 285 1194 287
rect 1138 283 1139 285
rect 1141 283 1142 285
rect 1174 284 1194 285
rect 1138 280 1142 283
rect 1118 276 1142 280
rect 1118 272 1122 276
rect 1164 280 1168 282
rect 1164 278 1165 280
rect 1167 278 1168 280
rect 1117 270 1122 272
rect 1117 268 1118 270
rect 1120 268 1122 270
rect 1126 271 1142 272
rect 1126 269 1128 271
rect 1130 269 1142 271
rect 1126 268 1142 269
rect 1117 266 1122 268
rect 1118 264 1122 266
rect 1118 261 1134 264
rect 1118 260 1131 261
rect 1130 259 1131 260
rect 1133 259 1134 261
rect 1130 254 1134 259
rect 1130 252 1131 254
rect 1133 252 1134 254
rect 1130 250 1134 252
rect 1138 262 1142 268
rect 1164 272 1168 278
rect 1157 268 1168 272
rect 1190 280 1194 284
rect 1205 281 1206 283
rect 1190 276 1202 280
rect 1198 271 1202 276
rect 1198 269 1199 271
rect 1201 269 1202 271
rect 1157 262 1161 268
rect 1138 261 1161 262
rect 1138 259 1157 261
rect 1159 259 1161 261
rect 1138 258 1161 259
rect 1073 245 1074 247
rect 1076 245 1077 247
rect 1073 243 1077 245
rect 1082 249 1088 250
rect 1082 247 1084 249
rect 1086 247 1088 249
rect 1138 247 1142 258
rect 1198 257 1202 269
rect 1185 254 1202 257
rect 1185 252 1186 254
rect 1188 253 1202 254
rect 1188 252 1189 253
rect 1082 238 1088 247
rect 1109 246 1142 247
rect 1109 244 1111 246
rect 1113 244 1142 246
rect 1109 243 1142 244
rect 1146 247 1150 249
rect 1146 245 1147 247
rect 1149 245 1150 247
rect 1146 240 1150 245
rect 1174 247 1180 248
rect 1174 245 1176 247
rect 1178 245 1180 247
rect 1146 238 1147 240
rect 1149 238 1150 240
rect 1174 238 1180 245
rect 1185 247 1189 252
rect 1185 245 1186 247
rect 1188 245 1189 247
rect 1185 243 1189 245
rect 1194 249 1200 250
rect 1194 247 1196 249
rect 1198 247 1200 249
rect 1194 238 1200 247
rect 12 220 14 222
rect 16 220 18 222
rect 12 219 18 220
rect 20 215 37 216
rect 20 213 33 215
rect 35 213 37 215
rect 20 212 37 213
rect 51 213 57 222
rect 5 201 6 212
rect 20 208 24 212
rect 51 211 53 213
rect 55 211 57 213
rect 51 210 57 211
rect 62 215 66 217
rect 62 213 63 215
rect 65 213 66 215
rect 9 204 24 208
rect 9 191 13 204
rect 62 208 66 213
rect 71 215 77 222
rect 101 220 102 222
rect 104 220 105 222
rect 71 213 73 215
rect 75 213 77 215
rect 71 212 77 213
rect 101 215 105 220
rect 101 213 102 215
rect 104 213 105 215
rect 101 211 105 213
rect 109 216 142 217
rect 109 214 138 216
rect 140 214 142 216
rect 109 213 142 214
rect 156 213 162 222
rect 62 207 63 208
rect 49 206 63 207
rect 65 206 66 208
rect 49 203 66 206
rect 28 195 34 196
rect 9 189 10 191
rect 12 189 13 191
rect 9 183 13 189
rect 9 182 27 183
rect 9 180 23 182
rect 25 180 27 182
rect 9 179 27 180
rect 49 191 53 203
rect 109 202 113 213
rect 156 211 158 213
rect 160 211 162 213
rect 156 210 162 211
rect 167 215 171 217
rect 167 213 168 215
rect 170 213 171 215
rect 90 201 113 202
rect 90 199 92 201
rect 94 199 113 201
rect 90 198 113 199
rect 90 192 94 198
rect 49 189 50 191
rect 52 189 53 191
rect 49 184 53 189
rect 49 180 61 184
rect 45 177 46 179
rect 57 176 61 180
rect 83 188 94 192
rect 83 182 87 188
rect 109 192 113 198
rect 117 208 121 210
rect 117 206 118 208
rect 120 206 121 208
rect 117 201 121 206
rect 117 199 118 201
rect 120 200 121 201
rect 120 199 133 200
rect 117 196 133 199
rect 129 194 133 196
rect 129 192 134 194
rect 109 191 125 192
rect 109 189 121 191
rect 123 189 125 191
rect 109 188 125 189
rect 129 190 131 192
rect 133 190 134 192
rect 129 188 134 190
rect 83 180 84 182
rect 86 180 87 182
rect 83 178 87 180
rect 129 184 133 188
rect 109 180 133 184
rect 109 177 113 180
rect 57 175 77 176
rect 109 175 110 177
rect 112 175 113 177
rect 57 173 73 175
rect 75 173 77 175
rect 57 172 77 173
rect 96 174 102 175
rect 96 172 98 174
rect 100 172 102 174
rect 109 173 113 175
rect 167 208 171 213
rect 176 215 182 222
rect 206 220 207 222
rect 209 220 210 222
rect 176 213 178 215
rect 180 213 182 215
rect 176 212 182 213
rect 206 215 210 220
rect 262 220 264 222
rect 266 220 268 222
rect 262 219 268 220
rect 206 213 207 215
rect 209 213 210 215
rect 206 211 210 213
rect 214 216 247 217
rect 214 214 243 216
rect 245 214 247 216
rect 214 213 247 214
rect 167 207 168 208
rect 154 206 168 207
rect 170 206 171 208
rect 154 203 171 206
rect 154 191 158 203
rect 214 202 218 213
rect 270 215 287 216
rect 270 213 283 215
rect 285 213 287 215
rect 270 212 287 213
rect 301 213 307 222
rect 195 201 218 202
rect 195 199 197 201
rect 199 199 218 201
rect 195 198 218 199
rect 195 192 199 198
rect 154 189 155 191
rect 157 189 158 191
rect 154 184 158 189
rect 154 180 166 184
rect 150 177 151 179
rect 12 169 18 170
rect 12 167 14 169
rect 16 167 18 169
rect 12 166 18 167
rect 31 169 37 170
rect 31 167 33 169
rect 35 167 37 169
rect 31 166 37 167
rect 96 166 102 172
rect 162 176 166 180
rect 188 188 199 192
rect 188 182 192 188
rect 214 192 218 198
rect 222 208 226 210
rect 222 206 223 208
rect 225 206 226 208
rect 222 201 226 206
rect 222 199 223 201
rect 225 200 226 201
rect 225 199 238 200
rect 222 196 238 199
rect 234 194 238 196
rect 234 192 239 194
rect 214 191 230 192
rect 214 189 226 191
rect 228 189 230 191
rect 214 188 230 189
rect 234 190 236 192
rect 238 190 239 192
rect 234 188 239 190
rect 188 180 189 182
rect 191 180 192 182
rect 188 178 192 180
rect 234 184 238 188
rect 214 180 238 184
rect 214 177 218 180
rect 162 175 182 176
rect 214 175 215 177
rect 217 175 218 177
rect 255 201 256 212
rect 270 208 274 212
rect 301 211 303 213
rect 305 211 307 213
rect 301 210 307 211
rect 312 215 316 217
rect 312 213 313 215
rect 315 213 316 215
rect 259 204 274 208
rect 259 191 263 204
rect 312 208 316 213
rect 321 215 327 222
rect 351 220 352 222
rect 354 220 355 222
rect 321 213 323 215
rect 325 213 327 215
rect 321 212 327 213
rect 351 215 355 220
rect 351 213 352 215
rect 354 213 355 215
rect 351 211 355 213
rect 359 216 392 217
rect 359 214 388 216
rect 390 214 392 216
rect 359 213 392 214
rect 406 213 412 222
rect 312 207 313 208
rect 299 206 313 207
rect 315 206 316 208
rect 299 203 316 206
rect 278 195 284 196
rect 259 189 260 191
rect 262 189 263 191
rect 259 183 263 189
rect 259 182 277 183
rect 259 180 273 182
rect 275 180 277 182
rect 259 179 277 180
rect 162 173 178 175
rect 180 173 182 175
rect 162 172 182 173
rect 201 174 207 175
rect 201 172 203 174
rect 205 172 207 174
rect 214 173 218 175
rect 299 191 303 203
rect 359 202 363 213
rect 406 211 408 213
rect 410 211 412 213
rect 406 210 412 211
rect 417 215 421 217
rect 417 213 418 215
rect 420 213 421 215
rect 340 201 363 202
rect 340 199 342 201
rect 344 199 363 201
rect 340 198 363 199
rect 340 192 344 198
rect 299 189 300 191
rect 302 189 303 191
rect 299 184 303 189
rect 299 180 311 184
rect 295 177 296 179
rect 201 166 207 172
rect 307 176 311 180
rect 333 188 344 192
rect 333 182 337 188
rect 359 192 363 198
rect 367 208 371 210
rect 367 206 368 208
rect 370 206 371 208
rect 367 201 371 206
rect 367 199 368 201
rect 370 200 371 201
rect 370 199 383 200
rect 367 196 383 199
rect 379 194 383 196
rect 379 192 384 194
rect 359 191 375 192
rect 359 189 371 191
rect 373 189 375 191
rect 359 188 375 189
rect 379 190 381 192
rect 383 190 384 192
rect 379 188 384 190
rect 333 180 334 182
rect 336 180 337 182
rect 333 178 337 180
rect 379 184 383 188
rect 359 180 383 184
rect 359 177 363 180
rect 307 175 327 176
rect 359 175 360 177
rect 362 175 363 177
rect 307 173 323 175
rect 325 173 327 175
rect 307 172 327 173
rect 346 174 352 175
rect 346 172 348 174
rect 350 172 352 174
rect 359 173 363 175
rect 417 208 421 213
rect 426 215 432 222
rect 456 220 457 222
rect 459 220 460 222
rect 426 213 428 215
rect 430 213 432 215
rect 426 212 432 213
rect 456 215 460 220
rect 512 220 514 222
rect 516 220 518 222
rect 512 219 518 220
rect 456 213 457 215
rect 459 213 460 215
rect 456 211 460 213
rect 464 216 497 217
rect 464 214 493 216
rect 495 214 497 216
rect 464 213 497 214
rect 417 207 418 208
rect 404 206 418 207
rect 420 206 421 208
rect 404 203 421 206
rect 404 191 408 203
rect 464 202 468 213
rect 520 215 537 216
rect 520 213 533 215
rect 535 213 537 215
rect 520 212 537 213
rect 551 213 557 222
rect 445 201 468 202
rect 445 199 447 201
rect 449 199 468 201
rect 445 198 468 199
rect 445 192 449 198
rect 404 189 405 191
rect 407 189 408 191
rect 404 184 408 189
rect 404 180 416 184
rect 400 177 401 179
rect 262 169 268 170
rect 262 167 264 169
rect 266 167 268 169
rect 262 166 268 167
rect 281 169 287 170
rect 281 167 283 169
rect 285 167 287 169
rect 281 166 287 167
rect 346 166 352 172
rect 412 176 416 180
rect 438 188 449 192
rect 438 182 442 188
rect 464 192 468 198
rect 472 208 476 210
rect 472 206 473 208
rect 475 206 476 208
rect 472 201 476 206
rect 472 199 473 201
rect 475 200 476 201
rect 475 199 488 200
rect 472 196 488 199
rect 484 194 488 196
rect 484 192 489 194
rect 464 191 480 192
rect 464 189 476 191
rect 478 189 480 191
rect 464 188 480 189
rect 484 190 486 192
rect 488 190 489 192
rect 484 188 489 190
rect 438 180 439 182
rect 441 180 442 182
rect 438 178 442 180
rect 484 184 488 188
rect 464 180 488 184
rect 464 177 468 180
rect 412 175 432 176
rect 464 175 465 177
rect 467 175 468 177
rect 505 201 506 212
rect 520 208 524 212
rect 551 211 553 213
rect 555 211 557 213
rect 551 210 557 211
rect 562 215 566 217
rect 562 213 563 215
rect 565 213 566 215
rect 509 204 524 208
rect 509 191 513 204
rect 562 208 566 213
rect 571 215 577 222
rect 601 220 602 222
rect 604 220 605 222
rect 571 213 573 215
rect 575 213 577 215
rect 571 212 577 213
rect 601 215 605 220
rect 601 213 602 215
rect 604 213 605 215
rect 601 211 605 213
rect 609 216 642 217
rect 609 214 638 216
rect 640 214 642 216
rect 609 213 642 214
rect 656 213 662 222
rect 562 207 563 208
rect 549 206 563 207
rect 565 206 566 208
rect 549 203 566 206
rect 528 195 534 196
rect 509 189 510 191
rect 512 189 513 191
rect 509 183 513 189
rect 509 182 527 183
rect 509 180 523 182
rect 525 180 527 182
rect 509 179 527 180
rect 412 173 428 175
rect 430 173 432 175
rect 412 172 432 173
rect 451 174 457 175
rect 451 172 453 174
rect 455 172 457 174
rect 464 173 468 175
rect 549 191 553 203
rect 609 202 613 213
rect 656 211 658 213
rect 660 211 662 213
rect 656 210 662 211
rect 667 215 671 217
rect 667 213 668 215
rect 670 213 671 215
rect 590 201 613 202
rect 590 199 592 201
rect 594 199 613 201
rect 590 198 613 199
rect 590 192 594 198
rect 549 189 550 191
rect 552 189 553 191
rect 549 184 553 189
rect 549 180 561 184
rect 545 177 546 179
rect 451 166 457 172
rect 557 176 561 180
rect 583 188 594 192
rect 583 182 587 188
rect 609 192 613 198
rect 617 208 621 210
rect 617 206 618 208
rect 620 206 621 208
rect 617 201 621 206
rect 617 199 618 201
rect 620 200 621 201
rect 620 199 633 200
rect 617 196 633 199
rect 629 194 633 196
rect 629 192 634 194
rect 609 191 625 192
rect 609 189 621 191
rect 623 189 625 191
rect 609 188 625 189
rect 629 190 631 192
rect 633 190 634 192
rect 629 188 634 190
rect 583 180 584 182
rect 586 180 587 182
rect 583 178 587 180
rect 629 184 633 188
rect 609 180 633 184
rect 609 177 613 180
rect 557 175 577 176
rect 609 175 610 177
rect 612 175 613 177
rect 557 173 573 175
rect 575 173 577 175
rect 557 172 577 173
rect 596 174 602 175
rect 596 172 598 174
rect 600 172 602 174
rect 609 173 613 175
rect 667 208 671 213
rect 676 215 682 222
rect 706 220 707 222
rect 709 220 710 222
rect 676 213 678 215
rect 680 213 682 215
rect 676 212 682 213
rect 706 215 710 220
rect 762 220 764 222
rect 766 220 768 222
rect 762 219 768 220
rect 706 213 707 215
rect 709 213 710 215
rect 706 211 710 213
rect 714 216 747 217
rect 714 214 743 216
rect 745 214 747 216
rect 714 213 747 214
rect 667 207 668 208
rect 654 206 668 207
rect 670 206 671 208
rect 654 203 671 206
rect 654 191 658 203
rect 714 202 718 213
rect 770 215 787 216
rect 770 213 783 215
rect 785 213 787 215
rect 770 212 787 213
rect 801 213 807 222
rect 695 201 718 202
rect 695 199 697 201
rect 699 199 718 201
rect 695 198 718 199
rect 695 192 699 198
rect 654 189 655 191
rect 657 189 658 191
rect 654 184 658 189
rect 654 180 666 184
rect 650 177 651 179
rect 512 169 518 170
rect 512 167 514 169
rect 516 167 518 169
rect 512 166 518 167
rect 531 169 537 170
rect 531 167 533 169
rect 535 167 537 169
rect 531 166 537 167
rect 596 166 602 172
rect 662 176 666 180
rect 688 188 699 192
rect 688 182 692 188
rect 714 192 718 198
rect 722 208 726 210
rect 722 206 723 208
rect 725 206 726 208
rect 722 201 726 206
rect 722 199 723 201
rect 725 200 726 201
rect 725 199 738 200
rect 722 196 738 199
rect 734 194 738 196
rect 734 192 739 194
rect 714 191 730 192
rect 714 189 726 191
rect 728 189 730 191
rect 714 188 730 189
rect 734 190 736 192
rect 738 190 739 192
rect 734 188 739 190
rect 688 180 689 182
rect 691 180 692 182
rect 688 178 692 180
rect 734 184 738 188
rect 714 180 738 184
rect 714 177 718 180
rect 662 175 682 176
rect 714 175 715 177
rect 717 175 718 177
rect 755 201 756 212
rect 770 208 774 212
rect 801 211 803 213
rect 805 211 807 213
rect 801 210 807 211
rect 812 215 816 217
rect 812 213 813 215
rect 815 213 816 215
rect 759 204 774 208
rect 759 191 763 204
rect 812 208 816 213
rect 821 215 827 222
rect 851 220 852 222
rect 854 220 855 222
rect 821 213 823 215
rect 825 213 827 215
rect 821 212 827 213
rect 851 215 855 220
rect 851 213 852 215
rect 854 213 855 215
rect 851 211 855 213
rect 859 216 892 217
rect 859 214 888 216
rect 890 214 892 216
rect 859 213 892 214
rect 906 213 912 222
rect 812 207 813 208
rect 799 206 813 207
rect 815 206 816 208
rect 799 203 816 206
rect 778 195 784 196
rect 759 189 760 191
rect 762 189 763 191
rect 759 183 763 189
rect 759 182 777 183
rect 759 180 773 182
rect 775 180 777 182
rect 759 179 777 180
rect 662 173 678 175
rect 680 173 682 175
rect 662 172 682 173
rect 701 174 707 175
rect 701 172 703 174
rect 705 172 707 174
rect 714 173 718 175
rect 799 191 803 203
rect 859 202 863 213
rect 906 211 908 213
rect 910 211 912 213
rect 906 210 912 211
rect 917 215 921 217
rect 917 213 918 215
rect 920 213 921 215
rect 840 201 863 202
rect 840 199 842 201
rect 844 199 863 201
rect 840 198 863 199
rect 840 192 844 198
rect 799 189 800 191
rect 802 189 803 191
rect 799 184 803 189
rect 799 180 811 184
rect 795 177 796 179
rect 701 166 707 172
rect 807 176 811 180
rect 833 188 844 192
rect 833 182 837 188
rect 859 192 863 198
rect 867 208 871 210
rect 867 206 868 208
rect 870 206 871 208
rect 867 201 871 206
rect 867 199 868 201
rect 870 200 871 201
rect 870 199 883 200
rect 867 196 883 199
rect 879 194 883 196
rect 879 192 884 194
rect 859 191 875 192
rect 859 189 871 191
rect 873 189 875 191
rect 859 188 875 189
rect 879 190 881 192
rect 883 190 884 192
rect 879 188 884 190
rect 833 180 834 182
rect 836 180 837 182
rect 833 178 837 180
rect 879 184 883 188
rect 859 180 883 184
rect 859 177 863 180
rect 807 175 827 176
rect 859 175 860 177
rect 862 175 863 177
rect 807 173 823 175
rect 825 173 827 175
rect 807 172 827 173
rect 846 174 852 175
rect 846 172 848 174
rect 850 172 852 174
rect 859 173 863 175
rect 917 208 921 213
rect 926 215 932 222
rect 956 220 957 222
rect 959 220 960 222
rect 926 213 928 215
rect 930 213 932 215
rect 926 212 932 213
rect 956 215 960 220
rect 956 213 957 215
rect 959 213 960 215
rect 956 211 960 213
rect 964 216 997 217
rect 964 214 993 216
rect 995 214 997 216
rect 964 213 997 214
rect 1032 213 1038 222
rect 917 207 918 208
rect 904 206 918 207
rect 920 206 921 208
rect 904 203 921 206
rect 904 191 908 203
rect 964 202 968 213
rect 1032 211 1034 213
rect 1036 211 1038 213
rect 1032 210 1038 211
rect 1043 215 1047 217
rect 1043 213 1044 215
rect 1046 213 1047 215
rect 945 201 968 202
rect 945 199 947 201
rect 949 199 968 201
rect 945 198 968 199
rect 945 192 949 198
rect 904 189 905 191
rect 907 189 908 191
rect 904 184 908 189
rect 904 180 916 184
rect 900 177 901 179
rect 762 169 768 170
rect 762 167 764 169
rect 766 167 768 169
rect 762 166 768 167
rect 781 169 787 170
rect 781 167 783 169
rect 785 167 787 169
rect 781 166 787 167
rect 846 166 852 172
rect 912 176 916 180
rect 938 188 949 192
rect 938 182 942 188
rect 964 192 968 198
rect 972 208 976 210
rect 972 206 973 208
rect 975 206 976 208
rect 972 201 976 206
rect 972 199 973 201
rect 975 200 976 201
rect 975 199 988 200
rect 972 196 988 199
rect 984 194 988 196
rect 984 192 989 194
rect 964 191 980 192
rect 964 189 976 191
rect 978 189 980 191
rect 964 188 980 189
rect 984 190 986 192
rect 988 190 989 192
rect 984 188 989 190
rect 938 180 939 182
rect 941 180 942 182
rect 938 178 942 180
rect 984 184 988 188
rect 964 180 988 184
rect 964 177 968 180
rect 912 175 932 176
rect 964 175 965 177
rect 967 175 968 177
rect 912 173 928 175
rect 930 173 932 175
rect 912 172 932 173
rect 951 174 957 175
rect 951 172 953 174
rect 955 172 957 174
rect 964 173 968 175
rect 1043 208 1047 213
rect 1052 215 1058 222
rect 1052 213 1054 215
rect 1056 213 1058 215
rect 1052 212 1058 213
rect 1062 215 1068 222
rect 1062 213 1064 215
rect 1066 213 1068 215
rect 1062 212 1068 213
rect 1073 215 1077 217
rect 1073 213 1074 215
rect 1076 213 1077 215
rect 1043 207 1044 208
rect 1030 206 1044 207
rect 1046 206 1047 208
rect 1030 203 1047 206
rect 1030 191 1034 203
rect 1073 208 1077 213
rect 1082 213 1088 222
rect 1082 211 1084 213
rect 1086 211 1088 213
rect 1082 210 1088 211
rect 1112 213 1118 222
rect 1112 211 1114 213
rect 1116 211 1118 213
rect 1112 210 1118 211
rect 1123 215 1127 217
rect 1123 213 1124 215
rect 1126 213 1127 215
rect 1073 206 1074 208
rect 1076 207 1077 208
rect 1076 206 1090 207
rect 1073 203 1090 206
rect 1030 189 1031 191
rect 1033 189 1034 191
rect 1030 184 1034 189
rect 1030 180 1042 184
rect 1026 177 1027 179
rect 951 166 957 172
rect 1038 176 1042 180
rect 1086 191 1090 203
rect 1086 189 1087 191
rect 1089 189 1090 191
rect 1086 184 1090 189
rect 1078 180 1090 184
rect 1078 176 1082 180
rect 1093 177 1094 179
rect 1038 175 1058 176
rect 1038 173 1054 175
rect 1056 173 1058 175
rect 1038 172 1058 173
rect 1062 175 1082 176
rect 1062 173 1064 175
rect 1066 173 1082 175
rect 1062 172 1082 173
rect 1123 208 1127 213
rect 1132 215 1138 222
rect 1162 220 1163 222
rect 1165 220 1166 222
rect 1132 213 1134 215
rect 1136 213 1138 215
rect 1132 212 1138 213
rect 1162 215 1166 220
rect 1162 213 1163 215
rect 1165 213 1166 215
rect 1162 211 1166 213
rect 1170 216 1203 217
rect 1170 214 1199 216
rect 1201 214 1203 216
rect 1170 213 1203 214
rect 1123 207 1124 208
rect 1110 206 1124 207
rect 1126 206 1127 208
rect 1110 203 1127 206
rect 1110 191 1114 203
rect 1170 202 1174 213
rect 1151 201 1174 202
rect 1151 199 1153 201
rect 1155 199 1174 201
rect 1151 198 1174 199
rect 1151 192 1155 198
rect 1110 189 1111 191
rect 1113 189 1114 191
rect 1110 184 1114 189
rect 1110 180 1122 184
rect 1106 177 1107 179
rect 1118 176 1122 180
rect 1144 188 1155 192
rect 1144 182 1148 188
rect 1170 192 1174 198
rect 1178 208 1182 210
rect 1178 206 1179 208
rect 1181 206 1182 208
rect 1178 201 1182 206
rect 1178 199 1179 201
rect 1181 200 1182 201
rect 1181 199 1194 200
rect 1178 196 1194 199
rect 1190 194 1194 196
rect 1190 192 1195 194
rect 1170 191 1186 192
rect 1170 189 1182 191
rect 1184 189 1186 191
rect 1170 188 1186 189
rect 1190 190 1192 192
rect 1194 190 1195 192
rect 1190 188 1195 190
rect 1144 180 1145 182
rect 1147 180 1148 182
rect 1144 178 1148 180
rect 1190 184 1194 188
rect 1170 180 1194 184
rect 1170 177 1174 180
rect 1118 175 1138 176
rect 1170 175 1171 177
rect 1173 175 1174 177
rect 1118 173 1134 175
rect 1136 173 1138 175
rect 1118 172 1138 173
rect 1157 174 1163 175
rect 1157 172 1159 174
rect 1161 172 1163 174
rect 1170 173 1174 175
rect 1157 166 1163 172
rect 155 135 161 141
rect 226 140 232 141
rect 226 138 228 140
rect 230 138 232 140
rect 226 137 232 138
rect 245 140 251 141
rect 245 138 247 140
rect 249 138 251 140
rect 245 137 251 138
rect 116 134 136 135
rect 116 132 132 134
rect 134 132 136 134
rect 155 133 157 135
rect 159 133 161 135
rect 155 132 161 133
rect 168 132 172 134
rect 116 131 136 132
rect 104 128 105 130
rect 116 127 120 131
rect 168 130 169 132
rect 171 130 172 132
rect 108 123 120 127
rect 108 118 112 123
rect 108 116 109 118
rect 111 116 112 118
rect 108 104 112 116
rect 142 127 146 129
rect 142 125 143 127
rect 145 125 146 127
rect 142 119 146 125
rect 168 127 172 130
rect 168 123 192 127
rect 142 115 153 119
rect 149 109 153 115
rect 188 119 192 123
rect 168 118 184 119
rect 168 116 180 118
rect 182 116 184 118
rect 168 115 184 116
rect 188 117 193 119
rect 188 115 190 117
rect 192 115 193 117
rect 168 109 172 115
rect 188 113 193 115
rect 310 135 316 141
rect 271 134 291 135
rect 271 132 287 134
rect 289 132 291 134
rect 310 133 312 135
rect 314 133 316 135
rect 310 132 316 133
rect 323 132 327 134
rect 271 131 291 132
rect 188 111 192 113
rect 149 108 172 109
rect 149 106 151 108
rect 153 106 172 108
rect 149 105 172 106
rect 108 101 125 104
rect 108 100 122 101
rect 121 99 122 100
rect 124 99 125 101
rect 110 96 116 97
rect 110 94 112 96
rect 114 94 116 96
rect 110 85 116 94
rect 121 94 125 99
rect 121 92 122 94
rect 124 92 125 94
rect 121 90 125 92
rect 130 94 136 95
rect 130 92 132 94
rect 134 92 136 94
rect 130 85 136 92
rect 160 94 164 96
rect 160 92 161 94
rect 163 92 164 94
rect 160 87 164 92
rect 168 94 172 105
rect 176 108 192 111
rect 176 106 177 108
rect 179 107 192 108
rect 179 106 180 107
rect 176 101 180 106
rect 176 99 177 101
rect 179 99 180 101
rect 176 97 180 99
rect 223 127 241 128
rect 223 125 237 127
rect 239 125 241 127
rect 223 124 241 125
rect 223 118 227 124
rect 259 128 260 130
rect 271 127 275 131
rect 323 130 324 132
rect 326 130 327 132
rect 223 116 224 118
rect 226 116 227 118
rect 219 95 220 106
rect 223 103 227 116
rect 242 111 248 112
rect 223 99 238 103
rect 234 95 238 99
rect 263 123 275 127
rect 263 118 267 123
rect 263 116 264 118
rect 266 116 267 118
rect 263 104 267 116
rect 297 127 301 129
rect 297 125 298 127
rect 300 125 301 127
rect 297 119 301 125
rect 323 127 327 130
rect 323 123 347 127
rect 297 115 308 119
rect 304 109 308 115
rect 343 119 347 123
rect 323 118 339 119
rect 323 116 335 118
rect 337 116 339 118
rect 323 115 339 116
rect 343 117 348 119
rect 343 115 345 117
rect 347 115 348 117
rect 323 109 327 115
rect 343 113 348 115
rect 343 111 347 113
rect 304 108 327 109
rect 304 106 306 108
rect 308 106 327 108
rect 304 105 327 106
rect 263 101 280 104
rect 263 100 277 101
rect 276 99 277 100
rect 279 99 280 101
rect 265 96 271 97
rect 168 93 201 94
rect 168 91 197 93
rect 199 91 201 93
rect 168 90 201 91
rect 234 94 251 95
rect 234 92 247 94
rect 249 92 251 94
rect 234 91 251 92
rect 265 94 267 96
rect 269 94 271 96
rect 160 85 161 87
rect 163 85 164 87
rect 226 87 232 88
rect 226 85 228 87
rect 230 85 232 87
rect 265 85 271 94
rect 276 94 280 99
rect 276 92 277 94
rect 279 92 280 94
rect 276 90 280 92
rect 285 94 291 95
rect 285 92 287 94
rect 289 92 291 94
rect 285 85 291 92
rect 315 94 319 96
rect 315 92 316 94
rect 318 92 319 94
rect 315 87 319 92
rect 323 94 327 105
rect 331 108 347 111
rect 331 106 332 108
rect 334 107 347 108
rect 334 106 335 107
rect 331 101 335 106
rect 331 99 332 101
rect 334 99 335 101
rect 331 97 335 99
rect 415 135 421 141
rect 476 140 482 141
rect 476 138 478 140
rect 480 138 482 140
rect 476 137 482 138
rect 495 140 501 141
rect 495 138 497 140
rect 499 138 501 140
rect 495 137 501 138
rect 376 134 396 135
rect 376 132 392 134
rect 394 132 396 134
rect 415 133 417 135
rect 419 133 421 135
rect 415 132 421 133
rect 428 132 432 134
rect 376 131 396 132
rect 364 128 365 130
rect 376 127 380 131
rect 428 130 429 132
rect 431 130 432 132
rect 368 123 380 127
rect 368 118 372 123
rect 368 116 369 118
rect 371 116 372 118
rect 368 104 372 116
rect 402 127 406 129
rect 402 125 403 127
rect 405 125 406 127
rect 402 119 406 125
rect 428 127 432 130
rect 428 123 452 127
rect 402 115 413 119
rect 409 109 413 115
rect 448 119 452 123
rect 428 118 444 119
rect 428 116 440 118
rect 442 116 444 118
rect 428 115 444 116
rect 448 117 453 119
rect 448 115 450 117
rect 452 115 453 117
rect 428 109 432 115
rect 448 113 453 115
rect 448 111 452 113
rect 409 108 432 109
rect 409 106 411 108
rect 413 106 432 108
rect 409 105 432 106
rect 368 101 385 104
rect 368 100 382 101
rect 381 99 382 100
rect 384 99 385 101
rect 370 96 376 97
rect 370 94 372 96
rect 374 94 376 96
rect 323 93 356 94
rect 323 91 352 93
rect 354 91 356 93
rect 323 90 356 91
rect 315 85 316 87
rect 318 85 319 87
rect 370 85 376 94
rect 381 94 385 99
rect 381 92 382 94
rect 384 92 385 94
rect 381 90 385 92
rect 390 94 396 95
rect 390 92 392 94
rect 394 92 396 94
rect 390 85 396 92
rect 420 94 424 96
rect 420 92 421 94
rect 423 92 424 94
rect 420 87 424 92
rect 428 94 432 105
rect 436 108 452 111
rect 436 106 437 108
rect 439 107 452 108
rect 439 106 440 107
rect 436 101 440 106
rect 560 135 566 141
rect 521 134 541 135
rect 521 132 537 134
rect 539 132 541 134
rect 560 133 562 135
rect 564 133 566 135
rect 560 132 566 133
rect 573 132 577 134
rect 521 131 541 132
rect 436 99 437 101
rect 439 99 440 101
rect 436 97 440 99
rect 473 127 491 128
rect 473 125 487 127
rect 489 125 491 127
rect 473 124 491 125
rect 473 118 477 124
rect 509 128 510 130
rect 521 127 525 131
rect 573 130 574 132
rect 576 130 577 132
rect 473 116 474 118
rect 476 116 477 118
rect 469 95 470 106
rect 473 103 477 116
rect 492 111 498 112
rect 473 99 488 103
rect 484 95 488 99
rect 513 123 525 127
rect 513 118 517 123
rect 513 116 514 118
rect 516 116 517 118
rect 513 104 517 116
rect 547 127 551 129
rect 547 125 548 127
rect 550 125 551 127
rect 547 119 551 125
rect 573 127 577 130
rect 573 123 597 127
rect 547 115 558 119
rect 554 109 558 115
rect 593 119 597 123
rect 573 118 589 119
rect 573 116 585 118
rect 587 116 589 118
rect 573 115 589 116
rect 593 117 598 119
rect 593 115 595 117
rect 597 115 598 117
rect 573 109 577 115
rect 593 113 598 115
rect 593 111 597 113
rect 554 108 577 109
rect 554 106 556 108
rect 558 106 577 108
rect 554 105 577 106
rect 513 101 530 104
rect 513 100 527 101
rect 526 99 527 100
rect 529 99 530 101
rect 515 96 521 97
rect 428 93 461 94
rect 428 91 457 93
rect 459 91 461 93
rect 428 90 461 91
rect 484 94 501 95
rect 484 92 497 94
rect 499 92 501 94
rect 484 91 501 92
rect 515 94 517 96
rect 519 94 521 96
rect 420 85 421 87
rect 423 85 424 87
rect 476 87 482 88
rect 476 85 478 87
rect 480 85 482 87
rect 515 85 521 94
rect 526 94 530 99
rect 526 92 527 94
rect 529 92 530 94
rect 526 90 530 92
rect 535 94 541 95
rect 535 92 537 94
rect 539 92 541 94
rect 535 85 541 92
rect 565 94 569 96
rect 565 92 566 94
rect 568 92 569 94
rect 565 87 569 92
rect 573 94 577 105
rect 581 108 597 111
rect 581 106 582 108
rect 584 107 597 108
rect 584 106 585 107
rect 581 101 585 106
rect 581 99 582 101
rect 584 99 585 101
rect 581 97 585 99
rect 665 135 671 141
rect 726 140 732 141
rect 726 138 728 140
rect 730 138 732 140
rect 726 137 732 138
rect 745 140 751 141
rect 745 138 747 140
rect 749 138 751 140
rect 745 137 751 138
rect 626 134 646 135
rect 626 132 642 134
rect 644 132 646 134
rect 665 133 667 135
rect 669 133 671 135
rect 665 132 671 133
rect 678 132 682 134
rect 626 131 646 132
rect 614 128 615 130
rect 626 127 630 131
rect 678 130 679 132
rect 681 130 682 132
rect 618 123 630 127
rect 618 118 622 123
rect 618 116 619 118
rect 621 116 622 118
rect 618 104 622 116
rect 652 127 656 129
rect 652 125 653 127
rect 655 125 656 127
rect 652 119 656 125
rect 678 127 682 130
rect 678 123 702 127
rect 652 115 663 119
rect 659 109 663 115
rect 698 119 702 123
rect 678 118 694 119
rect 678 116 690 118
rect 692 116 694 118
rect 678 115 694 116
rect 698 117 703 119
rect 698 115 700 117
rect 702 115 703 117
rect 678 109 682 115
rect 698 113 703 115
rect 698 111 702 113
rect 659 108 682 109
rect 659 106 661 108
rect 663 106 682 108
rect 659 105 682 106
rect 618 101 635 104
rect 618 100 632 101
rect 631 99 632 100
rect 634 99 635 101
rect 620 96 626 97
rect 620 94 622 96
rect 624 94 626 96
rect 573 93 606 94
rect 573 91 602 93
rect 604 91 606 93
rect 573 90 606 91
rect 565 85 566 87
rect 568 85 569 87
rect 620 85 626 94
rect 631 94 635 99
rect 631 92 632 94
rect 634 92 635 94
rect 631 90 635 92
rect 640 94 646 95
rect 640 92 642 94
rect 644 92 646 94
rect 640 85 646 92
rect 670 94 674 96
rect 670 92 671 94
rect 673 92 674 94
rect 670 87 674 92
rect 678 94 682 105
rect 686 108 702 111
rect 686 106 687 108
rect 689 107 702 108
rect 689 106 690 107
rect 686 101 690 106
rect 810 135 816 141
rect 771 134 791 135
rect 771 132 787 134
rect 789 132 791 134
rect 810 133 812 135
rect 814 133 816 135
rect 810 132 816 133
rect 823 132 827 134
rect 771 131 791 132
rect 686 99 687 101
rect 689 99 690 101
rect 686 97 690 99
rect 723 127 741 128
rect 723 125 737 127
rect 739 125 741 127
rect 723 124 741 125
rect 723 118 727 124
rect 759 128 760 130
rect 771 127 775 131
rect 823 130 824 132
rect 826 130 827 132
rect 723 116 724 118
rect 726 116 727 118
rect 719 95 720 106
rect 723 103 727 116
rect 742 111 748 112
rect 723 99 738 103
rect 734 95 738 99
rect 763 123 775 127
rect 763 118 767 123
rect 763 116 764 118
rect 766 116 767 118
rect 763 104 767 116
rect 797 127 801 129
rect 797 125 798 127
rect 800 125 801 127
rect 797 119 801 125
rect 823 127 827 130
rect 823 123 847 127
rect 797 115 808 119
rect 804 109 808 115
rect 843 119 847 123
rect 823 118 839 119
rect 823 116 835 118
rect 837 116 839 118
rect 823 115 839 116
rect 843 117 848 119
rect 843 115 845 117
rect 847 115 848 117
rect 823 109 827 115
rect 843 113 848 115
rect 843 111 847 113
rect 804 108 827 109
rect 804 106 806 108
rect 808 106 827 108
rect 804 105 827 106
rect 763 101 780 104
rect 763 100 777 101
rect 776 99 777 100
rect 779 99 780 101
rect 765 96 771 97
rect 678 93 711 94
rect 678 91 707 93
rect 709 91 711 93
rect 678 90 711 91
rect 734 94 751 95
rect 734 92 747 94
rect 749 92 751 94
rect 734 91 751 92
rect 765 94 767 96
rect 769 94 771 96
rect 670 85 671 87
rect 673 85 674 87
rect 726 87 732 88
rect 726 85 728 87
rect 730 85 732 87
rect 765 85 771 94
rect 776 94 780 99
rect 776 92 777 94
rect 779 92 780 94
rect 776 90 780 92
rect 785 94 791 95
rect 785 92 787 94
rect 789 92 791 94
rect 785 85 791 92
rect 815 94 819 96
rect 815 92 816 94
rect 818 92 819 94
rect 815 87 819 92
rect 823 94 827 105
rect 831 108 847 111
rect 831 106 832 108
rect 834 107 847 108
rect 834 106 835 107
rect 831 101 835 106
rect 831 99 832 101
rect 834 99 835 101
rect 831 97 835 99
rect 915 135 921 141
rect 976 140 982 141
rect 976 138 978 140
rect 980 138 982 140
rect 976 137 982 138
rect 995 140 1001 141
rect 995 138 997 140
rect 999 138 1001 140
rect 995 137 1001 138
rect 876 134 896 135
rect 876 132 892 134
rect 894 132 896 134
rect 915 133 917 135
rect 919 133 921 135
rect 915 132 921 133
rect 928 132 932 134
rect 876 131 896 132
rect 864 128 865 130
rect 876 127 880 131
rect 928 130 929 132
rect 931 130 932 132
rect 868 123 880 127
rect 868 118 872 123
rect 868 116 869 118
rect 871 116 872 118
rect 868 104 872 116
rect 902 127 906 129
rect 902 125 903 127
rect 905 125 906 127
rect 902 119 906 125
rect 928 127 932 130
rect 928 123 952 127
rect 902 115 913 119
rect 909 109 913 115
rect 948 119 952 123
rect 928 118 944 119
rect 928 116 940 118
rect 942 116 944 118
rect 928 115 944 116
rect 948 117 953 119
rect 948 115 950 117
rect 952 115 953 117
rect 928 109 932 115
rect 948 113 953 115
rect 948 111 952 113
rect 909 108 932 109
rect 909 106 911 108
rect 913 106 932 108
rect 909 105 932 106
rect 868 101 885 104
rect 868 100 882 101
rect 881 99 882 100
rect 884 99 885 101
rect 870 96 876 97
rect 870 94 872 96
rect 874 94 876 96
rect 823 93 856 94
rect 823 91 852 93
rect 854 91 856 93
rect 823 90 856 91
rect 815 85 816 87
rect 818 85 819 87
rect 870 85 876 94
rect 881 94 885 99
rect 881 92 882 94
rect 884 92 885 94
rect 881 90 885 92
rect 890 94 896 95
rect 890 92 892 94
rect 894 92 896 94
rect 890 85 896 92
rect 920 94 924 96
rect 920 92 921 94
rect 923 92 924 94
rect 920 87 924 92
rect 928 94 932 105
rect 936 108 952 111
rect 936 106 937 108
rect 939 107 952 108
rect 939 106 940 107
rect 936 101 940 106
rect 1060 135 1066 141
rect 1021 134 1041 135
rect 1021 132 1037 134
rect 1039 132 1041 134
rect 1060 133 1062 135
rect 1064 133 1066 135
rect 1060 132 1066 133
rect 1073 132 1077 134
rect 1021 131 1041 132
rect 936 99 937 101
rect 939 99 940 101
rect 936 97 940 99
rect 973 127 991 128
rect 973 125 987 127
rect 989 125 991 127
rect 973 124 991 125
rect 973 118 977 124
rect 1009 128 1010 130
rect 1021 127 1025 131
rect 1073 130 1074 132
rect 1076 130 1077 132
rect 973 116 974 118
rect 976 116 977 118
rect 969 95 970 106
rect 973 103 977 116
rect 992 111 998 112
rect 973 99 988 103
rect 984 95 988 99
rect 1013 123 1025 127
rect 1013 118 1017 123
rect 1013 116 1014 118
rect 1016 116 1017 118
rect 1013 104 1017 116
rect 1047 127 1051 129
rect 1047 125 1048 127
rect 1050 125 1051 127
rect 1047 119 1051 125
rect 1073 127 1077 130
rect 1073 123 1097 127
rect 1047 115 1058 119
rect 1054 109 1058 115
rect 1093 119 1097 123
rect 1073 118 1089 119
rect 1073 116 1085 118
rect 1087 116 1089 118
rect 1073 115 1089 116
rect 1093 117 1098 119
rect 1093 115 1095 117
rect 1097 115 1098 117
rect 1073 109 1077 115
rect 1093 113 1098 115
rect 1093 111 1097 113
rect 1054 108 1077 109
rect 1054 106 1056 108
rect 1058 106 1077 108
rect 1054 105 1077 106
rect 1013 101 1030 104
rect 1013 100 1027 101
rect 1026 99 1027 100
rect 1029 99 1030 101
rect 1015 96 1021 97
rect 928 93 961 94
rect 928 91 957 93
rect 959 91 961 93
rect 928 90 961 91
rect 984 94 1001 95
rect 984 92 997 94
rect 999 92 1001 94
rect 984 91 1001 92
rect 1015 94 1017 96
rect 1019 94 1021 96
rect 920 85 921 87
rect 923 85 924 87
rect 976 87 982 88
rect 976 85 978 87
rect 980 85 982 87
rect 1015 85 1021 94
rect 1026 94 1030 99
rect 1026 92 1027 94
rect 1029 92 1030 94
rect 1026 90 1030 92
rect 1035 94 1041 95
rect 1035 92 1037 94
rect 1039 92 1041 94
rect 1035 85 1041 92
rect 1065 94 1069 96
rect 1065 92 1066 94
rect 1068 92 1069 94
rect 1065 87 1069 92
rect 1073 94 1077 105
rect 1081 108 1097 111
rect 1081 106 1082 108
rect 1084 107 1097 108
rect 1084 106 1085 107
rect 1081 101 1085 106
rect 1081 99 1082 101
rect 1084 99 1085 101
rect 1081 97 1085 99
rect 1165 135 1171 141
rect 1126 134 1146 135
rect 1126 132 1142 134
rect 1144 132 1146 134
rect 1165 133 1167 135
rect 1169 133 1171 135
rect 1165 132 1171 133
rect 1178 132 1182 134
rect 1126 131 1146 132
rect 1114 128 1115 130
rect 1126 127 1130 131
rect 1178 130 1179 132
rect 1181 130 1182 132
rect 1118 123 1130 127
rect 1118 118 1122 123
rect 1118 116 1119 118
rect 1121 116 1122 118
rect 1118 104 1122 116
rect 1152 127 1156 129
rect 1152 125 1153 127
rect 1155 125 1156 127
rect 1152 119 1156 125
rect 1178 127 1182 130
rect 1178 123 1202 127
rect 1152 115 1163 119
rect 1159 109 1163 115
rect 1198 119 1202 123
rect 1178 118 1194 119
rect 1178 116 1190 118
rect 1192 116 1194 118
rect 1178 115 1194 116
rect 1198 117 1203 119
rect 1198 115 1200 117
rect 1202 115 1203 117
rect 1178 109 1182 115
rect 1198 113 1203 115
rect 1198 111 1202 113
rect 1159 108 1182 109
rect 1159 106 1161 108
rect 1163 106 1182 108
rect 1159 105 1182 106
rect 1118 101 1135 104
rect 1118 100 1132 101
rect 1131 99 1132 100
rect 1134 99 1135 101
rect 1120 96 1126 97
rect 1120 94 1122 96
rect 1124 94 1126 96
rect 1073 93 1106 94
rect 1073 91 1102 93
rect 1104 91 1106 93
rect 1073 90 1106 91
rect 1065 85 1066 87
rect 1068 85 1069 87
rect 1120 85 1126 94
rect 1131 94 1135 99
rect 1131 92 1132 94
rect 1134 92 1135 94
rect 1131 90 1135 92
rect 1140 94 1146 95
rect 1140 92 1142 94
rect 1144 92 1146 94
rect 1140 85 1146 92
rect 1170 94 1174 96
rect 1170 92 1171 94
rect 1173 92 1174 94
rect 1170 87 1174 92
rect 1178 94 1182 105
rect 1186 108 1202 111
rect 1186 106 1187 108
rect 1189 107 1202 108
rect 1189 106 1190 107
rect 1186 101 1190 106
rect 1186 99 1187 101
rect 1189 99 1190 101
rect 1186 97 1190 99
rect 1178 93 1211 94
rect 1178 91 1207 93
rect 1209 91 1211 93
rect 1178 90 1211 91
rect 1170 85 1171 87
rect 1173 85 1174 87
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 26 62 43 63
rect 26 60 39 62
rect 41 60 43 62
rect 26 59 43 60
rect 57 60 63 69
rect 11 48 12 59
rect 26 55 30 59
rect 57 58 59 60
rect 61 58 63 60
rect 57 57 63 58
rect 68 62 72 64
rect 68 60 69 62
rect 71 60 72 62
rect 15 51 30 55
rect 15 38 19 51
rect 68 55 72 60
rect 77 62 83 69
rect 107 67 108 69
rect 110 67 111 69
rect 77 60 79 62
rect 81 60 83 62
rect 77 59 83 60
rect 107 62 111 67
rect 107 60 108 62
rect 110 60 111 62
rect 107 58 111 60
rect 115 63 148 64
rect 115 61 144 63
rect 146 61 148 63
rect 115 60 148 61
rect 162 60 168 69
rect 68 54 69 55
rect 55 53 69 54
rect 71 53 72 55
rect 55 50 72 53
rect 34 42 40 43
rect 15 36 16 38
rect 18 36 19 38
rect 15 30 19 36
rect 15 29 33 30
rect 15 27 29 29
rect 31 27 33 29
rect 15 26 33 27
rect 55 38 59 50
rect 115 49 119 60
rect 162 58 164 60
rect 166 58 168 60
rect 162 57 168 58
rect 173 62 177 64
rect 173 60 174 62
rect 176 60 177 62
rect 96 48 119 49
rect 96 46 98 48
rect 100 46 119 48
rect 96 45 119 46
rect 96 39 100 45
rect 55 36 56 38
rect 58 36 59 38
rect 55 31 59 36
rect 55 27 67 31
rect 51 24 52 26
rect 63 23 67 27
rect 89 35 100 39
rect 89 29 93 35
rect 115 39 119 45
rect 123 55 127 57
rect 123 53 124 55
rect 126 53 127 55
rect 123 48 127 53
rect 123 46 124 48
rect 126 47 127 48
rect 126 46 139 47
rect 123 43 139 46
rect 135 41 139 43
rect 135 39 140 41
rect 115 38 131 39
rect 115 36 127 38
rect 129 36 131 38
rect 115 35 131 36
rect 135 37 137 39
rect 139 37 140 39
rect 135 35 140 37
rect 89 27 90 29
rect 92 27 93 29
rect 89 25 93 27
rect 135 31 139 35
rect 115 27 139 31
rect 115 24 119 27
rect 63 22 83 23
rect 115 22 116 24
rect 118 22 119 24
rect 63 20 79 22
rect 81 20 83 22
rect 63 19 83 20
rect 102 21 108 22
rect 102 19 104 21
rect 106 19 108 21
rect 115 20 119 22
rect 173 55 177 60
rect 182 62 188 69
rect 212 67 213 69
rect 215 67 216 69
rect 182 60 184 62
rect 186 60 188 62
rect 182 59 188 60
rect 212 62 216 67
rect 268 67 270 69
rect 272 67 274 69
rect 268 66 274 67
rect 212 60 213 62
rect 215 60 216 62
rect 212 58 216 60
rect 220 63 253 64
rect 220 61 249 63
rect 251 61 253 63
rect 220 60 253 61
rect 173 54 174 55
rect 160 53 174 54
rect 176 53 177 55
rect 160 50 177 53
rect 160 38 164 50
rect 220 49 224 60
rect 276 62 293 63
rect 276 60 289 62
rect 291 60 293 62
rect 276 59 293 60
rect 307 60 313 69
rect 201 48 224 49
rect 201 46 203 48
rect 205 46 224 48
rect 201 45 224 46
rect 201 39 205 45
rect 160 36 161 38
rect 163 36 164 38
rect 160 31 164 36
rect 160 27 172 31
rect 156 24 157 26
rect 18 16 24 17
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 37 16 43 17
rect 37 14 39 16
rect 41 14 43 16
rect 37 13 43 14
rect 102 13 108 19
rect 168 23 172 27
rect 194 35 205 39
rect 194 29 198 35
rect 220 39 224 45
rect 228 55 232 57
rect 228 53 229 55
rect 231 53 232 55
rect 228 48 232 53
rect 228 46 229 48
rect 231 47 232 48
rect 231 46 244 47
rect 228 43 244 46
rect 240 41 244 43
rect 240 39 245 41
rect 220 38 236 39
rect 220 36 232 38
rect 234 36 236 38
rect 220 35 236 36
rect 240 37 242 39
rect 244 37 245 39
rect 240 35 245 37
rect 194 27 195 29
rect 197 27 198 29
rect 194 25 198 27
rect 240 31 244 35
rect 220 27 244 31
rect 220 24 224 27
rect 168 22 188 23
rect 220 22 221 24
rect 223 22 224 24
rect 261 48 262 59
rect 276 55 280 59
rect 307 58 309 60
rect 311 58 313 60
rect 307 57 313 58
rect 318 62 322 64
rect 318 60 319 62
rect 321 60 322 62
rect 265 51 280 55
rect 265 38 269 51
rect 318 55 322 60
rect 327 62 333 69
rect 357 67 358 69
rect 360 67 361 69
rect 327 60 329 62
rect 331 60 333 62
rect 327 59 333 60
rect 357 62 361 67
rect 357 60 358 62
rect 360 60 361 62
rect 357 58 361 60
rect 365 63 398 64
rect 365 61 394 63
rect 396 61 398 63
rect 365 60 398 61
rect 412 60 418 69
rect 318 54 319 55
rect 305 53 319 54
rect 321 53 322 55
rect 305 50 322 53
rect 284 42 290 43
rect 265 36 266 38
rect 268 36 269 38
rect 265 30 269 36
rect 265 29 283 30
rect 265 27 279 29
rect 281 27 283 29
rect 265 26 283 27
rect 168 20 184 22
rect 186 20 188 22
rect 168 19 188 20
rect 207 21 213 22
rect 207 19 209 21
rect 211 19 213 21
rect 220 20 224 22
rect 305 38 309 50
rect 365 49 369 60
rect 412 58 414 60
rect 416 58 418 60
rect 412 57 418 58
rect 423 62 427 64
rect 423 60 424 62
rect 426 60 427 62
rect 346 48 369 49
rect 346 46 348 48
rect 350 46 369 48
rect 346 45 369 46
rect 346 39 350 45
rect 305 36 306 38
rect 308 36 309 38
rect 305 31 309 36
rect 305 27 317 31
rect 301 24 302 26
rect 207 13 213 19
rect 313 23 317 27
rect 339 35 350 39
rect 339 29 343 35
rect 365 39 369 45
rect 373 55 377 57
rect 373 53 374 55
rect 376 53 377 55
rect 373 48 377 53
rect 373 46 374 48
rect 376 47 377 48
rect 376 46 389 47
rect 373 43 389 46
rect 385 41 389 43
rect 385 39 390 41
rect 365 38 381 39
rect 365 36 377 38
rect 379 36 381 38
rect 365 35 381 36
rect 385 37 387 39
rect 389 37 390 39
rect 385 35 390 37
rect 339 27 340 29
rect 342 27 343 29
rect 339 25 343 27
rect 385 31 389 35
rect 365 27 389 31
rect 365 24 369 27
rect 313 22 333 23
rect 365 22 366 24
rect 368 22 369 24
rect 313 20 329 22
rect 331 20 333 22
rect 313 19 333 20
rect 352 21 358 22
rect 352 19 354 21
rect 356 19 358 21
rect 365 20 369 22
rect 423 55 427 60
rect 432 62 438 69
rect 462 67 463 69
rect 465 67 466 69
rect 432 60 434 62
rect 436 60 438 62
rect 432 59 438 60
rect 462 62 466 67
rect 518 67 520 69
rect 522 67 524 69
rect 518 66 524 67
rect 462 60 463 62
rect 465 60 466 62
rect 462 58 466 60
rect 470 63 503 64
rect 470 61 499 63
rect 501 61 503 63
rect 470 60 503 61
rect 423 54 424 55
rect 410 53 424 54
rect 426 53 427 55
rect 410 50 427 53
rect 410 38 414 50
rect 470 49 474 60
rect 526 62 543 63
rect 526 60 539 62
rect 541 60 543 62
rect 526 59 543 60
rect 557 60 563 69
rect 451 48 474 49
rect 451 46 453 48
rect 455 46 474 48
rect 451 45 474 46
rect 451 39 455 45
rect 410 36 411 38
rect 413 36 414 38
rect 410 31 414 36
rect 410 27 422 31
rect 406 24 407 26
rect 268 16 274 17
rect 268 14 270 16
rect 272 14 274 16
rect 268 13 274 14
rect 287 16 293 17
rect 287 14 289 16
rect 291 14 293 16
rect 287 13 293 14
rect 352 13 358 19
rect 418 23 422 27
rect 444 35 455 39
rect 444 29 448 35
rect 470 39 474 45
rect 478 55 482 57
rect 478 53 479 55
rect 481 53 482 55
rect 478 48 482 53
rect 478 46 479 48
rect 481 47 482 48
rect 481 46 494 47
rect 478 43 494 46
rect 490 41 494 43
rect 490 39 495 41
rect 470 38 486 39
rect 470 36 482 38
rect 484 36 486 38
rect 470 35 486 36
rect 490 37 492 39
rect 494 37 495 39
rect 490 35 495 37
rect 444 27 445 29
rect 447 27 448 29
rect 444 25 448 27
rect 490 31 494 35
rect 470 27 494 31
rect 470 24 474 27
rect 418 22 438 23
rect 470 22 471 24
rect 473 22 474 24
rect 511 48 512 59
rect 526 55 530 59
rect 557 58 559 60
rect 561 58 563 60
rect 557 57 563 58
rect 568 62 572 64
rect 568 60 569 62
rect 571 60 572 62
rect 515 51 530 55
rect 515 38 519 51
rect 568 55 572 60
rect 577 62 583 69
rect 607 67 608 69
rect 610 67 611 69
rect 577 60 579 62
rect 581 60 583 62
rect 577 59 583 60
rect 607 62 611 67
rect 607 60 608 62
rect 610 60 611 62
rect 607 58 611 60
rect 615 63 648 64
rect 615 61 644 63
rect 646 61 648 63
rect 615 60 648 61
rect 662 60 668 69
rect 568 54 569 55
rect 555 53 569 54
rect 571 53 572 55
rect 555 50 572 53
rect 534 42 540 43
rect 515 36 516 38
rect 518 36 519 38
rect 515 30 519 36
rect 515 29 533 30
rect 515 27 529 29
rect 531 27 533 29
rect 515 26 533 27
rect 418 20 434 22
rect 436 20 438 22
rect 418 19 438 20
rect 457 21 463 22
rect 457 19 459 21
rect 461 19 463 21
rect 470 20 474 22
rect 555 38 559 50
rect 615 49 619 60
rect 662 58 664 60
rect 666 58 668 60
rect 662 57 668 58
rect 673 62 677 64
rect 673 60 674 62
rect 676 60 677 62
rect 596 48 619 49
rect 596 46 598 48
rect 600 46 619 48
rect 596 45 619 46
rect 596 39 600 45
rect 555 36 556 38
rect 558 36 559 38
rect 555 31 559 36
rect 555 27 567 31
rect 551 24 552 26
rect 457 13 463 19
rect 563 23 567 27
rect 589 35 600 39
rect 589 29 593 35
rect 615 39 619 45
rect 623 55 627 57
rect 623 53 624 55
rect 626 53 627 55
rect 623 48 627 53
rect 623 46 624 48
rect 626 47 627 48
rect 626 46 639 47
rect 623 43 639 46
rect 635 41 639 43
rect 635 39 640 41
rect 615 38 631 39
rect 615 36 627 38
rect 629 36 631 38
rect 615 35 631 36
rect 635 37 637 39
rect 639 37 640 39
rect 635 35 640 37
rect 589 27 590 29
rect 592 27 593 29
rect 589 25 593 27
rect 635 31 639 35
rect 615 27 639 31
rect 615 24 619 27
rect 563 22 583 23
rect 615 22 616 24
rect 618 22 619 24
rect 563 20 579 22
rect 581 20 583 22
rect 563 19 583 20
rect 602 21 608 22
rect 602 19 604 21
rect 606 19 608 21
rect 615 20 619 22
rect 673 55 677 60
rect 682 62 688 69
rect 712 67 713 69
rect 715 67 716 69
rect 682 60 684 62
rect 686 60 688 62
rect 682 59 688 60
rect 712 62 716 67
rect 768 67 770 69
rect 772 67 774 69
rect 768 66 774 67
rect 712 60 713 62
rect 715 60 716 62
rect 712 58 716 60
rect 720 63 753 64
rect 720 61 749 63
rect 751 61 753 63
rect 720 60 753 61
rect 673 54 674 55
rect 660 53 674 54
rect 676 53 677 55
rect 660 50 677 53
rect 660 38 664 50
rect 720 49 724 60
rect 776 62 793 63
rect 776 60 789 62
rect 791 60 793 62
rect 776 59 793 60
rect 807 60 813 69
rect 701 48 724 49
rect 701 46 703 48
rect 705 46 724 48
rect 701 45 724 46
rect 701 39 705 45
rect 660 36 661 38
rect 663 36 664 38
rect 660 31 664 36
rect 660 27 672 31
rect 656 24 657 26
rect 518 16 524 17
rect 518 14 520 16
rect 522 14 524 16
rect 518 13 524 14
rect 537 16 543 17
rect 537 14 539 16
rect 541 14 543 16
rect 537 13 543 14
rect 602 13 608 19
rect 668 23 672 27
rect 694 35 705 39
rect 694 29 698 35
rect 720 39 724 45
rect 728 55 732 57
rect 728 53 729 55
rect 731 53 732 55
rect 728 48 732 53
rect 728 46 729 48
rect 731 47 732 48
rect 731 46 744 47
rect 728 43 744 46
rect 740 41 744 43
rect 740 39 745 41
rect 720 38 736 39
rect 720 36 732 38
rect 734 36 736 38
rect 720 35 736 36
rect 740 37 742 39
rect 744 37 745 39
rect 740 35 745 37
rect 694 27 695 29
rect 697 27 698 29
rect 694 25 698 27
rect 740 31 744 35
rect 720 27 744 31
rect 720 24 724 27
rect 668 22 688 23
rect 720 22 721 24
rect 723 22 724 24
rect 761 48 762 59
rect 776 55 780 59
rect 807 58 809 60
rect 811 58 813 60
rect 807 57 813 58
rect 818 62 822 64
rect 818 60 819 62
rect 821 60 822 62
rect 765 51 780 55
rect 765 38 769 51
rect 818 55 822 60
rect 827 62 833 69
rect 857 67 858 69
rect 860 67 861 69
rect 827 60 829 62
rect 831 60 833 62
rect 827 59 833 60
rect 857 62 861 67
rect 857 60 858 62
rect 860 60 861 62
rect 857 58 861 60
rect 865 63 898 64
rect 865 61 894 63
rect 896 61 898 63
rect 865 60 898 61
rect 912 60 918 69
rect 818 54 819 55
rect 805 53 819 54
rect 821 53 822 55
rect 805 50 822 53
rect 784 42 790 43
rect 765 36 766 38
rect 768 36 769 38
rect 765 30 769 36
rect 765 29 783 30
rect 765 27 779 29
rect 781 27 783 29
rect 765 26 783 27
rect 668 20 684 22
rect 686 20 688 22
rect 668 19 688 20
rect 707 21 713 22
rect 707 19 709 21
rect 711 19 713 21
rect 720 20 724 22
rect 805 38 809 50
rect 865 49 869 60
rect 912 58 914 60
rect 916 58 918 60
rect 912 57 918 58
rect 923 62 927 64
rect 923 60 924 62
rect 926 60 927 62
rect 846 48 869 49
rect 846 46 848 48
rect 850 46 869 48
rect 846 45 869 46
rect 846 39 850 45
rect 805 36 806 38
rect 808 36 809 38
rect 805 31 809 36
rect 805 27 817 31
rect 801 24 802 26
rect 707 13 713 19
rect 813 23 817 27
rect 839 35 850 39
rect 839 29 843 35
rect 865 39 869 45
rect 873 55 877 57
rect 873 53 874 55
rect 876 53 877 55
rect 873 48 877 53
rect 873 46 874 48
rect 876 47 877 48
rect 876 46 889 47
rect 873 43 889 46
rect 885 41 889 43
rect 885 39 890 41
rect 865 38 881 39
rect 865 36 877 38
rect 879 36 881 38
rect 865 35 881 36
rect 885 37 887 39
rect 889 37 890 39
rect 885 35 890 37
rect 839 27 840 29
rect 842 27 843 29
rect 839 25 843 27
rect 885 31 889 35
rect 865 27 889 31
rect 865 24 869 27
rect 813 22 833 23
rect 865 22 866 24
rect 868 22 869 24
rect 813 20 829 22
rect 831 20 833 22
rect 813 19 833 20
rect 852 21 858 22
rect 852 19 854 21
rect 856 19 858 21
rect 865 20 869 22
rect 923 55 927 60
rect 932 62 938 69
rect 962 67 963 69
rect 965 67 966 69
rect 932 60 934 62
rect 936 60 938 62
rect 932 59 938 60
rect 962 62 966 67
rect 962 60 963 62
rect 965 60 966 62
rect 962 58 966 60
rect 970 63 1003 64
rect 970 61 999 63
rect 1001 61 1003 63
rect 970 60 1003 61
rect 923 54 924 55
rect 910 53 924 54
rect 926 53 927 55
rect 910 50 927 53
rect 910 38 914 50
rect 970 49 974 60
rect 951 48 974 49
rect 951 46 953 48
rect 955 46 974 48
rect 951 45 974 46
rect 951 39 955 45
rect 910 36 911 38
rect 913 36 914 38
rect 910 31 914 36
rect 910 27 922 31
rect 906 24 907 26
rect 768 16 774 17
rect 768 14 770 16
rect 772 14 774 16
rect 768 13 774 14
rect 787 16 793 17
rect 787 14 789 16
rect 791 14 793 16
rect 787 13 793 14
rect 852 13 858 19
rect 918 23 922 27
rect 944 35 955 39
rect 944 29 948 35
rect 970 39 974 45
rect 978 55 982 57
rect 978 53 979 55
rect 981 53 982 55
rect 978 48 982 53
rect 978 46 979 48
rect 981 47 982 48
rect 981 46 994 47
rect 978 43 994 46
rect 990 41 994 43
rect 990 39 995 41
rect 970 38 986 39
rect 970 36 982 38
rect 984 36 986 38
rect 970 35 986 36
rect 990 37 992 39
rect 994 37 995 39
rect 990 35 995 37
rect 944 27 945 29
rect 947 27 948 29
rect 944 25 948 27
rect 990 31 994 35
rect 970 27 994 31
rect 970 24 974 27
rect 918 22 938 23
rect 970 22 971 24
rect 973 22 974 24
rect 918 20 934 22
rect 936 20 938 22
rect 918 19 938 20
rect 957 21 963 22
rect 957 19 959 21
rect 961 19 963 21
rect 970 20 974 22
rect 957 13 963 19
<< via1 >>
rect 32 385 34 387
rect 47 394 49 396
rect 72 385 74 387
rect 15 369 17 371
rect 55 370 57 372
rect 86 371 88 373
rect 148 394 150 396
rect 175 394 177 396
rect 514 387 516 389
rect 199 382 201 384
rect 167 371 169 373
rect 529 396 531 398
rect 554 387 556 389
rect 497 371 499 373
rect 537 372 539 374
rect 568 373 570 375
rect 630 396 632 398
rect 657 396 659 398
rect 719 387 721 389
rect 681 384 683 386
rect 649 373 651 375
rect 734 396 736 398
rect 759 387 761 389
rect 702 371 704 373
rect 742 372 744 374
rect 773 373 775 375
rect 835 396 837 398
rect 862 396 864 398
rect 886 384 888 386
rect 854 373 856 375
rect 47 322 49 324
rect 55 313 57 315
rect 30 305 32 307
rect 72 305 74 307
rect 87 296 89 298
rect 143 329 145 331
rect 119 296 121 298
rect 146 296 148 298
rect 529 324 531 326
rect 537 315 539 317
rect 512 307 514 309
rect 554 307 556 309
rect 569 298 571 300
rect 625 331 627 333
rect 601 298 603 300
rect 628 298 630 300
rect 734 324 736 326
rect 742 315 744 317
rect 717 307 719 309
rect 759 307 761 309
rect 774 298 776 300
rect 830 331 832 333
rect 806 298 808 300
rect 833 298 835 300
rect 1040 269 1042 271
rect 1055 278 1057 280
rect 1080 269 1082 271
rect 1023 253 1025 255
rect 1063 254 1065 256
rect 1094 255 1096 257
rect 1156 278 1158 280
rect 1183 278 1185 280
rect 1207 266 1209 268
rect 1175 255 1177 257
rect 34 206 36 208
rect 3 180 5 182
rect 66 180 68 182
rect 93 180 95 182
rect 139 180 141 182
rect 148 206 150 208
rect 181 198 183 200
rect 171 180 173 182
rect 198 180 200 182
rect 284 206 286 208
rect 252 198 254 200
rect 316 180 318 182
rect 343 180 345 182
rect 389 180 391 182
rect 398 206 400 208
rect 433 198 435 200
rect 421 180 423 182
rect 448 180 450 182
rect 534 206 536 208
rect 502 198 504 200
rect 566 180 568 182
rect 593 180 595 182
rect 639 180 641 182
rect 648 206 650 208
rect 683 198 685 200
rect 671 180 673 182
rect 698 180 700 182
rect 784 206 786 208
rect 752 198 754 200
rect 816 180 818 182
rect 843 180 845 182
rect 889 180 891 182
rect 898 206 900 208
rect 921 180 923 182
rect 948 180 950 182
rect 1055 206 1057 208
rect 1063 197 1065 199
rect 1038 189 1040 191
rect 1080 189 1082 191
rect 1095 180 1097 182
rect 1151 213 1153 215
rect 1127 180 1129 182
rect 1154 180 1156 182
rect 1200 176 1202 178
rect 308 143 310 145
rect 558 142 560 144
rect 1147 143 1149 145
rect 125 125 127 127
rect 102 99 104 101
rect 116 116 118 118
rect 152 125 154 127
rect 143 108 145 110
rect 198 111 200 113
rect 217 125 219 127
rect 248 99 250 101
rect 280 125 282 127
rect 307 125 309 127
rect 353 125 355 127
rect 385 125 387 127
rect 362 99 364 101
rect 412 125 414 127
rect 395 107 397 109
rect 458 99 460 101
rect 466 107 468 109
rect 498 99 500 101
rect 530 125 532 127
rect 557 125 559 127
rect 603 125 605 127
rect 635 125 637 127
rect 612 99 614 101
rect 662 125 664 127
rect 647 107 649 109
rect 708 99 710 101
rect 716 107 718 109
rect 748 99 750 101
rect 780 125 782 127
rect 807 125 809 127
rect 853 125 855 127
rect 885 125 887 127
rect 862 99 864 101
rect 912 125 914 127
rect 897 107 899 109
rect 966 107 968 109
rect 998 99 1000 101
rect 1030 125 1032 127
rect 1057 125 1059 127
rect 1103 125 1105 127
rect 1135 125 1137 127
rect 1112 99 1114 101
rect 1162 125 1164 127
rect 1147 108 1149 110
rect 40 53 42 55
rect 72 27 74 29
rect 106 36 108 38
rect 99 27 101 29
rect 145 27 147 29
rect 154 53 156 55
rect 187 45 189 47
rect 177 27 179 29
rect 204 27 206 29
rect 290 53 292 55
rect 258 45 260 47
rect 322 27 324 29
rect 356 37 358 39
rect 349 27 351 29
rect 395 27 397 29
rect 404 53 406 55
rect 439 45 441 47
rect 427 27 429 29
rect 454 27 456 29
rect 540 53 542 55
rect 508 45 510 47
rect 572 27 574 29
rect 606 37 608 39
rect 599 27 601 29
rect 645 27 647 29
rect 654 53 656 55
rect 689 45 691 47
rect 677 27 679 29
rect 704 27 706 29
rect 790 53 792 55
rect 758 45 760 47
rect 822 27 824 29
rect 856 36 858 38
rect 849 27 851 29
rect 895 27 897 29
rect 904 53 906 55
rect 939 44 941 46
rect 927 27 929 29
rect 954 27 956 29
rect 939 9 941 11
<< via2 >>
rect 1103 188 1105 190
rect 1103 169 1105 171
rect 1147 133 1149 135
rect 1147 117 1149 119
rect 939 35 941 37
rect 939 19 941 21
<< labels >>
rlabel alu1 9 44 9 44 1 c2
rlabel alu1 98 61 98 61 1 p33
rlabel alu1 348 61 348 61 1 p32
rlabel alu1 598 61 598 61 1 p31
rlabel alu1 607 36 607 36 1 s13
rlabel alu1 848 61 848 61 1 p30
rlabel alu1 857 36 857 36 1 s12
rlabel alu1 1001 40 1001 40 1 r4
rlabel alu1 751 40 751 40 1 r5
rlabel alu1 501 40 501 40 1 r6
rlabel alu1 251 40 251 40 1 r7
rlabel alu1 357 36 357 36 1 sha
rlabel alu1 107 36 107 36 1 cha
rlabel alu1 285 9 285 9 1 Gnd
rlabel alu1 936 53 936 53 1 Gnd
rlabel alu1 1144 226 1144 226 1 Vdd
rlabel alu1 1120 226 1120 226 6 vdd
rlabel alu1 1142 161 1142 161 1 Vss
rlabel alu1 1040 162 1040 162 6 vss
rlabel alu1 1040 226 1040 226 6 vdd
rlabel alu1 1048 184 1048 184 1 a0
rlabel alu1 1056 206 1056 206 1 b0
rlabel alu1 1064 206 1064 206 1 b1
rlabel alu1 1072 185 1072 185 1 a1
rlabel alu1 1080 162 1080 162 4 vss
rlabel alu1 1080 226 1080 226 4 vdd
rlabel alu1 1170 299 1170 299 5 Vss
rlabel alu1 1192 234 1192 234 2 vdd
rlabel alu1 1168 234 1168 234 5 Vdd
rlabel alu1 1040 234 1040 234 2 vdd
rlabel alu1 1040 298 1040 298 2 vss
rlabel alu1 1080 298 1080 298 2 vss
rlabel alu1 1080 234 1080 234 2 vdd
rlabel alu1 1072 262 1072 262 1 b0
rlabel alu1 1072 274 1072 274 1 a1
rlabel alu1 1032 276 1032 276 1 a0
rlabel via1 1024 254 1024 254 1 b1
rlabel alu1 1024 190 1024 190 1 r0
rlabel alu1 1111 267 1111 267 1 r1
rlabel alu1 1201 193 1201 193 1 p02
rlabel alu1 1104 188 1104 188 1 p03
rlabel alu1 83 226 83 226 1 Vdd
rlabel alu1 59 226 59 226 6 vdd
rlabel alu1 81 161 81 161 1 Vss
rlabel alu1 188 226 188 226 1 Vdd
rlabel alu1 164 226 164 226 6 vdd
rlabel alu1 186 161 186 161 1 Vss
rlabel alu1 19 226 19 226 6 vdd
rlabel alu1 333 226 333 226 1 Vdd
rlabel alu1 309 226 309 226 6 vdd
rlabel alu1 331 161 331 161 1 Vss
rlabel alu1 438 226 438 226 1 Vdd
rlabel alu1 414 226 414 226 6 vdd
rlabel alu1 436 161 436 161 1 Vss
rlabel alu1 269 226 269 226 6 vdd
rlabel alu1 519 226 519 226 6 vdd
rlabel alu1 686 161 686 161 1 Vss
rlabel alu1 664 226 664 226 6 vdd
rlabel alu1 688 226 688 226 1 Vdd
rlabel alu1 581 161 581 161 1 Vss
rlabel alu1 559 226 559 226 6 vdd
rlabel alu1 583 226 583 226 1 Vdd
rlabel alu1 833 226 833 226 1 Vdd
rlabel alu1 809 226 809 226 6 vdd
rlabel alu1 831 161 831 161 1 Vss
rlabel alu1 938 226 938 226 1 Vdd
rlabel alu1 914 226 914 226 6 vdd
rlabel alu1 936 161 936 161 1 Vss
rlabel alu1 769 226 769 226 6 vdd
rlabel alu1 92 214 92 214 1 p23
rlabel alu1 101 189 101 189 1 p13
rlabel alu1 342 214 342 214 1 p22
rlabel alu1 351 189 351 189 1 p12
rlabel alu1 592 214 592 214 1 p21
rlabel alu1 601 189 601 189 1 p11
rlabel alu1 842 214 842 214 1 p20
rlabel alu1 851 189 851 189 1 p10
rlabel alu1 930 206 930 206 5 Vss
rlabel alu1 3 197 3 197 5 c0
rlabel alu1 245 193 245 193 5 s03
rlabel alu1 495 193 495 193 5 s02
rlabel alu1 745 193 745 193 5 s01
rlabel alu1 995 193 995 193 5 s00
rlabel alu1 618 344 618 344 1 Vdd
rlabel alu1 594 344 594 344 6 vdd
rlabel alu1 616 279 616 279 1 Vss
rlabel alu1 514 280 514 280 6 vss
rlabel alu1 514 344 514 344 6 vdd
rlabel alu1 554 280 554 280 4 vss
rlabel alu1 554 344 554 344 4 vdd
rlabel alu1 644 417 644 417 5 Vss
rlabel alu1 666 352 666 352 2 vdd
rlabel alu1 642 352 642 352 5 Vdd
rlabel alu1 514 352 514 352 2 vdd
rlabel alu1 514 416 514 416 2 vss
rlabel alu1 554 416 554 416 2 vss
rlabel alu1 554 352 554 352 2 vdd
rlabel alu1 711 394 711 394 1 a0
rlabel alu1 751 392 751 392 1 a1
rlabel alu1 759 352 759 352 2 vdd
rlabel alu1 759 416 759 416 2 vss
rlabel alu1 719 416 719 416 2 vss
rlabel alu1 719 352 719 352 2 vdd
rlabel alu1 847 352 847 352 5 Vdd
rlabel alu1 871 352 871 352 2 vdd
rlabel alu1 849 417 849 417 5 Vss
rlabel alu1 759 344 759 344 4 vdd
rlabel alu1 759 280 759 280 4 vss
rlabel alu1 751 303 751 303 1 a1
rlabel alu1 727 302 727 302 1 a0
rlabel alu1 719 344 719 344 6 vdd
rlabel alu1 719 280 719 280 6 vss
rlabel alu1 821 279 821 279 1 Vss
rlabel alu1 799 344 799 344 6 vdd
rlabel alu1 823 344 823 344 1 Vdd
rlabel alu1 783 306 783 306 1 p13
rlabel alu1 703 308 703 308 1 p10
rlabel alu1 880 311 880 311 1 p12
rlabel alu1 790 385 790 385 1 p11
rlabel alu1 498 308 498 308 1 p20
rlabel alu1 578 306 578 306 1 p23
rlabel alu1 675 311 675 311 1 p22
rlabel via1 735 324 735 324 1 b2
rlabel alu1 743 324 743 324 1 b3
rlabel alu1 751 380 751 380 1 b2
rlabel via1 703 372 703 372 1 b3
rlabel via1 498 372 498 372 1 b1
rlabel alu1 546 380 546 380 1 b0
rlabel via1 530 324 530 324 1 b0
rlabel alu1 538 324 538 324 1 b1
rlabel alu1 522 302 522 302 1 a2
rlabel alu1 546 303 546 303 1 a3
rlabel alu1 506 394 506 394 1 a2
rlabel alu1 546 392 546 392 1 a3
rlabel alu1 585 385 585 385 1 p21
rlabel alu1 1144 101 1144 101 1 Gnd
rlabel alu1 1209 114 1209 114 5 s10
rlabel alu1 959 114 959 114 5 s11
rlabel alu1 709 114 709 114 5 s12
rlabel alu1 459 114 459 114 5 s13
rlabel alu1 217 110 217 110 5 c1
rlabel alu1 306 93 306 93 5 s03
rlabel alu1 315 118 315 118 5 Vss
rlabel alu1 556 93 556 93 5 s02
rlabel alu1 565 118 565 118 5 Vss
rlabel alu1 806 93 806 93 5 s01
rlabel alu1 815 118 815 118 5 p03
rlabel alu1 1056 93 1056 93 5 s00
rlabel alu1 1065 118 1065 118 5 p02
rlabel alu1 983 81 983 81 8 vdd
rlabel alu1 1128 81 1128 81 8 vdd
rlabel alu1 1152 81 1152 81 5 Vdd
rlabel alu1 1023 81 1023 81 8 vdd
rlabel alu1 1047 81 1047 81 5 Vdd
rlabel alu1 797 81 797 81 5 Vdd
rlabel alu1 773 81 773 81 8 vdd
rlabel alu1 902 81 902 81 5 Vdd
rlabel alu1 878 81 878 81 8 vdd
rlabel alu1 733 81 733 81 8 vdd
rlabel alu1 483 81 483 81 8 vdd
rlabel alu1 628 81 628 81 8 vdd
rlabel alu1 652 81 652 81 5 Vdd
rlabel alu1 523 81 523 81 8 vdd
rlabel alu1 547 81 547 81 5 Vdd
rlabel alu1 233 81 233 81 8 vdd
rlabel alu1 378 81 378 81 8 vdd
rlabel alu1 402 81 402 81 5 Vdd
rlabel alu1 273 81 273 81 8 vdd
rlabel alu1 297 81 297 81 5 Vdd
rlabel alu1 140 146 140 146 1 Gnd
rlabel alu1 102 119 102 119 5 cha
rlabel alu1 151 93 151 93 5 c1
rlabel alu1 134 101 134 101 5 c1
rlabel alu1 160 118 160 118 5 c0
rlabel alu1 126 121 126 121 5 c0
rlabel alu1 199 114 199 114 5 sha
rlabel alu1 142 81 142 81 5 Vdd
rlabel alu1 136 342 136 342 1 Vdd
rlabel alu1 112 342 112 342 6 vdd
rlabel alu1 134 277 134 277 1 Vss
rlabel alu1 32 278 32 278 6 vss
rlabel alu1 32 342 32 342 6 vdd
rlabel alu1 72 278 72 278 4 vss
rlabel alu1 72 342 72 342 4 vdd
rlabel alu1 162 415 162 415 5 Vss
rlabel alu1 184 350 184 350 2 vdd
rlabel alu1 160 350 160 350 5 Vdd
rlabel alu1 32 350 32 350 2 vdd
rlabel alu1 32 414 32 414 2 vss
rlabel alu1 72 414 72 414 2 vss
rlabel alu1 72 350 72 350 2 vdd
rlabel alu1 40 300 40 300 1 a2
rlabel via1 48 322 48 322 1 b2
rlabel alu1 56 322 56 322 1 b3
rlabel alu1 64 301 64 301 1 a3
rlabel alu1 64 378 64 378 1 b2
rlabel alu1 64 390 64 390 1 a3
rlabel via1 16 370 16 370 1 b3
rlabel alu1 24 392 24 392 1 a2
rlabel alu1 16 306 16 306 1 p30
rlabel alu1 96 304 96 304 1 p33
rlabel alu1 193 309 193 309 1 p32
rlabel alu1 103 383 103 383 1 p31
<< end >>
