magic
tech scmos
timestamp 1608973495
<< ab >>
rect 5 5 85 77
rect 87 22 190 77
rect 87 13 100 22
rect 102 13 190 22
rect 87 5 190 13
rect 192 5 335 77
rect 337 5 440 77
rect 442 5 585 77
rect 587 5 690 77
rect 692 5 835 77
rect 837 34 940 77
rect 942 34 1005 77
rect 837 32 1005 34
rect 837 5 940 32
rect 942 5 1005 32
<< nwell >>
rect 0 37 1010 82
<< pwell >>
rect 0 0 1010 37
<< poly >>
rect 27 71 29 75
rect 34 71 36 75
rect 14 61 16 66
rect 103 71 105 75
rect 54 62 56 66
rect 64 64 66 69
rect 74 64 76 69
rect 14 40 16 43
rect 27 40 29 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 31 16 34
rect 24 31 26 34
rect 34 31 36 41
rect 54 40 56 44
rect 64 40 66 51
rect 74 48 76 51
rect 74 46 80 48
rect 74 44 76 46
rect 78 44 80 46
rect 74 42 80 44
rect 88 46 94 48
rect 88 44 90 46
rect 92 44 94 46
rect 139 71 141 75
rect 119 62 121 66
rect 129 62 131 66
rect 208 71 210 75
rect 159 62 161 66
rect 169 64 171 69
rect 179 64 181 69
rect 88 42 94 44
rect 54 38 60 40
rect 54 36 56 38
rect 58 36 60 38
rect 54 34 60 36
rect 64 38 70 40
rect 64 36 66 38
rect 68 36 70 38
rect 64 34 70 36
rect 54 29 56 34
rect 67 29 69 34
rect 74 29 76 42
rect 92 41 94 42
rect 103 41 105 44
rect 119 41 121 44
rect 92 39 105 41
rect 111 39 121 41
rect 129 40 131 44
rect 139 41 141 44
rect 95 31 97 39
rect 111 35 113 39
rect 104 33 113 35
rect 125 38 131 40
rect 125 36 127 38
rect 129 36 131 38
rect 125 34 131 36
rect 135 39 141 41
rect 135 37 137 39
rect 139 37 141 39
rect 135 35 141 37
rect 159 40 161 44
rect 169 40 171 51
rect 179 48 181 51
rect 179 46 185 48
rect 179 44 181 46
rect 183 44 185 46
rect 179 42 185 44
rect 193 46 199 48
rect 193 44 195 46
rect 197 44 199 46
rect 244 71 246 75
rect 224 62 226 66
rect 234 62 236 66
rect 277 71 279 75
rect 284 71 286 75
rect 264 61 266 66
rect 193 42 199 44
rect 159 38 165 40
rect 159 36 161 38
rect 163 36 165 38
rect 104 31 106 33
rect 108 31 113 33
rect 14 17 16 22
rect 24 20 26 25
rect 34 20 36 25
rect 54 16 56 20
rect 104 29 113 31
rect 129 31 131 34
rect 111 26 113 29
rect 121 26 123 30
rect 129 29 133 31
rect 131 26 133 29
rect 138 26 140 35
rect 159 34 165 36
rect 169 38 175 40
rect 169 36 171 38
rect 173 36 175 38
rect 169 34 175 36
rect 159 29 161 34
rect 172 29 174 34
rect 179 29 181 42
rect 197 41 199 42
rect 208 41 210 44
rect 224 41 226 44
rect 197 39 210 41
rect 216 39 226 41
rect 234 40 236 44
rect 244 41 246 44
rect 353 71 355 75
rect 304 62 306 66
rect 314 64 316 69
rect 324 64 326 69
rect 200 31 202 39
rect 216 35 218 39
rect 209 33 218 35
rect 230 38 236 40
rect 230 36 232 38
rect 234 36 236 38
rect 230 34 236 36
rect 240 39 246 41
rect 240 37 242 39
rect 244 37 246 39
rect 240 35 246 37
rect 264 40 266 43
rect 277 40 279 50
rect 284 47 286 50
rect 284 45 290 47
rect 284 43 286 45
rect 288 43 290 45
rect 284 41 290 43
rect 264 38 270 40
rect 264 36 266 38
rect 268 36 270 38
rect 209 31 211 33
rect 213 31 218 33
rect 95 19 97 22
rect 67 13 69 18
rect 74 13 76 18
rect 95 17 100 19
rect 98 9 100 17
rect 111 13 113 17
rect 121 9 123 17
rect 159 16 161 20
rect 209 29 218 31
rect 234 31 236 34
rect 216 26 218 29
rect 226 26 228 30
rect 234 29 238 31
rect 236 26 238 29
rect 243 26 245 35
rect 264 34 270 36
rect 274 38 280 40
rect 274 36 276 38
rect 278 36 280 38
rect 274 34 280 36
rect 264 31 266 34
rect 274 31 276 34
rect 284 31 286 41
rect 304 40 306 44
rect 314 40 316 51
rect 324 48 326 51
rect 324 46 330 48
rect 324 44 326 46
rect 328 44 330 46
rect 324 42 330 44
rect 338 46 344 48
rect 338 44 340 46
rect 342 44 344 46
rect 389 71 391 75
rect 369 62 371 66
rect 379 62 381 66
rect 458 71 460 75
rect 409 62 411 66
rect 419 64 421 69
rect 429 64 431 69
rect 338 42 344 44
rect 304 38 310 40
rect 304 36 306 38
rect 308 36 310 38
rect 304 34 310 36
rect 314 38 320 40
rect 314 36 316 38
rect 318 36 320 38
rect 314 34 320 36
rect 200 19 202 22
rect 131 9 133 14
rect 138 9 140 14
rect 98 7 123 9
rect 172 13 174 18
rect 179 13 181 18
rect 200 17 205 19
rect 203 9 205 17
rect 216 13 218 17
rect 226 9 228 17
rect 304 29 306 34
rect 317 29 319 34
rect 324 29 326 42
rect 342 41 344 42
rect 353 41 355 44
rect 369 41 371 44
rect 342 39 355 41
rect 361 39 371 41
rect 379 40 381 44
rect 389 41 391 44
rect 345 31 347 39
rect 361 35 363 39
rect 354 33 363 35
rect 375 38 381 40
rect 375 36 377 38
rect 379 36 381 38
rect 375 34 381 36
rect 385 39 391 41
rect 385 37 387 39
rect 389 37 391 39
rect 385 35 391 37
rect 409 40 411 44
rect 419 40 421 51
rect 429 48 431 51
rect 429 46 435 48
rect 429 44 431 46
rect 433 44 435 46
rect 429 42 435 44
rect 443 46 449 48
rect 443 44 445 46
rect 447 44 449 46
rect 494 71 496 75
rect 474 62 476 66
rect 484 62 486 66
rect 527 71 529 75
rect 534 71 536 75
rect 514 61 516 66
rect 443 42 449 44
rect 409 38 415 40
rect 409 36 411 38
rect 413 36 415 38
rect 354 31 356 33
rect 358 31 363 33
rect 264 17 266 22
rect 274 20 276 25
rect 284 20 286 25
rect 236 9 238 14
rect 243 9 245 14
rect 203 7 228 9
rect 304 16 306 20
rect 354 29 363 31
rect 379 31 381 34
rect 361 26 363 29
rect 371 26 373 30
rect 379 29 383 31
rect 381 26 383 29
rect 388 26 390 35
rect 409 34 415 36
rect 419 38 425 40
rect 419 36 421 38
rect 423 36 425 38
rect 419 34 425 36
rect 409 29 411 34
rect 422 29 424 34
rect 429 29 431 42
rect 447 41 449 42
rect 458 41 460 44
rect 474 41 476 44
rect 447 39 460 41
rect 466 39 476 41
rect 484 40 486 44
rect 494 41 496 44
rect 603 71 605 75
rect 554 62 556 66
rect 564 64 566 69
rect 574 64 576 69
rect 450 31 452 39
rect 466 35 468 39
rect 459 33 468 35
rect 480 38 486 40
rect 480 36 482 38
rect 484 36 486 38
rect 480 34 486 36
rect 490 39 496 41
rect 490 37 492 39
rect 494 37 496 39
rect 490 35 496 37
rect 514 40 516 43
rect 527 40 529 50
rect 534 47 536 50
rect 534 45 540 47
rect 534 43 536 45
rect 538 43 540 45
rect 534 41 540 43
rect 514 38 520 40
rect 514 36 516 38
rect 518 36 520 38
rect 459 31 461 33
rect 463 31 468 33
rect 345 19 347 22
rect 317 13 319 18
rect 324 13 326 18
rect 345 17 350 19
rect 348 9 350 17
rect 361 13 363 17
rect 371 9 373 17
rect 409 16 411 20
rect 459 29 468 31
rect 484 31 486 34
rect 466 26 468 29
rect 476 26 478 30
rect 484 29 488 31
rect 486 26 488 29
rect 493 26 495 35
rect 514 34 520 36
rect 524 38 530 40
rect 524 36 526 38
rect 528 36 530 38
rect 524 34 530 36
rect 514 31 516 34
rect 524 31 526 34
rect 534 31 536 41
rect 554 40 556 44
rect 564 40 566 51
rect 574 48 576 51
rect 574 46 580 48
rect 574 44 576 46
rect 578 44 580 46
rect 574 42 580 44
rect 588 46 594 48
rect 588 44 590 46
rect 592 44 594 46
rect 639 71 641 75
rect 619 62 621 66
rect 629 62 631 66
rect 708 71 710 75
rect 659 62 661 66
rect 669 64 671 69
rect 679 64 681 69
rect 588 42 594 44
rect 554 38 560 40
rect 554 36 556 38
rect 558 36 560 38
rect 554 34 560 36
rect 564 38 570 40
rect 564 36 566 38
rect 568 36 570 38
rect 564 34 570 36
rect 450 19 452 22
rect 381 9 383 14
rect 388 9 390 14
rect 348 7 373 9
rect 422 13 424 18
rect 429 13 431 18
rect 450 17 455 19
rect 453 9 455 17
rect 466 13 468 17
rect 476 9 478 17
rect 554 29 556 34
rect 567 29 569 34
rect 574 29 576 42
rect 592 41 594 42
rect 603 41 605 44
rect 619 41 621 44
rect 592 39 605 41
rect 611 39 621 41
rect 629 40 631 44
rect 639 41 641 44
rect 595 31 597 39
rect 611 35 613 39
rect 604 33 613 35
rect 625 38 631 40
rect 625 36 627 38
rect 629 36 631 38
rect 625 34 631 36
rect 635 39 641 41
rect 635 37 637 39
rect 639 37 641 39
rect 635 35 641 37
rect 659 40 661 44
rect 669 40 671 51
rect 679 48 681 51
rect 679 46 685 48
rect 679 44 681 46
rect 683 44 685 46
rect 679 42 685 44
rect 693 46 699 48
rect 693 44 695 46
rect 697 44 699 46
rect 744 71 746 75
rect 724 62 726 66
rect 734 62 736 66
rect 777 71 779 75
rect 784 71 786 75
rect 764 61 766 66
rect 693 42 699 44
rect 659 38 665 40
rect 659 36 661 38
rect 663 36 665 38
rect 604 31 606 33
rect 608 31 613 33
rect 514 17 516 22
rect 524 20 526 25
rect 534 20 536 25
rect 486 9 488 14
rect 493 9 495 14
rect 453 7 478 9
rect 554 16 556 20
rect 604 29 613 31
rect 629 31 631 34
rect 611 26 613 29
rect 621 26 623 30
rect 629 29 633 31
rect 631 26 633 29
rect 638 26 640 35
rect 659 34 665 36
rect 669 38 675 40
rect 669 36 671 38
rect 673 36 675 38
rect 669 34 675 36
rect 659 29 661 34
rect 672 29 674 34
rect 679 29 681 42
rect 697 41 699 42
rect 708 41 710 44
rect 724 41 726 44
rect 697 39 710 41
rect 716 39 726 41
rect 734 40 736 44
rect 744 41 746 44
rect 853 71 855 75
rect 804 62 806 66
rect 814 64 816 69
rect 824 64 826 69
rect 700 31 702 39
rect 716 35 718 39
rect 709 33 718 35
rect 730 38 736 40
rect 730 36 732 38
rect 734 36 736 38
rect 730 34 736 36
rect 740 39 746 41
rect 740 37 742 39
rect 744 37 746 39
rect 740 35 746 37
rect 764 40 766 43
rect 777 40 779 50
rect 784 47 786 50
rect 784 45 790 47
rect 784 43 786 45
rect 788 43 790 45
rect 784 41 790 43
rect 764 38 770 40
rect 764 36 766 38
rect 768 36 770 38
rect 709 31 711 33
rect 713 31 718 33
rect 595 19 597 22
rect 567 13 569 18
rect 574 13 576 18
rect 595 17 600 19
rect 598 9 600 17
rect 611 13 613 17
rect 621 9 623 17
rect 659 16 661 20
rect 709 29 718 31
rect 734 31 736 34
rect 716 26 718 29
rect 726 26 728 30
rect 734 29 738 31
rect 736 26 738 29
rect 743 26 745 35
rect 764 34 770 36
rect 774 38 780 40
rect 774 36 776 38
rect 778 36 780 38
rect 774 34 780 36
rect 764 31 766 34
rect 774 31 776 34
rect 784 31 786 41
rect 804 40 806 44
rect 814 40 816 51
rect 824 48 826 51
rect 824 46 830 48
rect 824 44 826 46
rect 828 44 830 46
rect 824 42 830 44
rect 838 46 844 48
rect 838 44 840 46
rect 842 44 844 46
rect 889 71 891 75
rect 869 62 871 66
rect 879 62 881 66
rect 958 71 960 75
rect 909 62 911 66
rect 919 64 921 69
rect 929 64 931 69
rect 838 42 844 44
rect 804 38 810 40
rect 804 36 806 38
rect 808 36 810 38
rect 804 34 810 36
rect 814 38 820 40
rect 814 36 816 38
rect 818 36 820 38
rect 814 34 820 36
rect 700 19 702 22
rect 631 9 633 14
rect 638 9 640 14
rect 598 7 623 9
rect 672 13 674 18
rect 679 13 681 18
rect 700 17 705 19
rect 703 9 705 17
rect 716 13 718 17
rect 726 9 728 17
rect 804 29 806 34
rect 817 29 819 34
rect 824 29 826 42
rect 842 41 844 42
rect 853 41 855 44
rect 869 41 871 44
rect 842 39 855 41
rect 861 39 871 41
rect 879 40 881 44
rect 889 41 891 44
rect 845 31 847 39
rect 861 35 863 39
rect 854 33 863 35
rect 875 38 881 40
rect 875 36 877 38
rect 879 36 881 38
rect 875 34 881 36
rect 885 39 891 41
rect 885 37 887 39
rect 889 37 891 39
rect 885 35 891 37
rect 909 40 911 44
rect 919 40 921 51
rect 929 48 931 51
rect 929 46 935 48
rect 929 44 931 46
rect 933 44 935 46
rect 929 42 935 44
rect 943 46 949 48
rect 943 44 945 46
rect 947 44 949 46
rect 994 71 996 75
rect 974 62 976 66
rect 984 62 986 66
rect 943 42 949 44
rect 909 38 915 40
rect 909 36 911 38
rect 913 36 915 38
rect 854 31 856 33
rect 858 31 863 33
rect 764 17 766 22
rect 774 20 776 25
rect 784 20 786 25
rect 736 9 738 14
rect 743 9 745 14
rect 703 7 728 9
rect 804 16 806 20
rect 854 29 863 31
rect 879 31 881 34
rect 861 26 863 29
rect 871 26 873 30
rect 879 29 883 31
rect 881 26 883 29
rect 888 26 890 35
rect 909 34 915 36
rect 919 38 925 40
rect 919 36 921 38
rect 923 36 925 38
rect 919 34 925 36
rect 909 29 911 34
rect 922 29 924 34
rect 929 29 931 42
rect 947 41 949 42
rect 958 41 960 44
rect 974 41 976 44
rect 947 39 960 41
rect 966 39 976 41
rect 984 40 986 44
rect 994 41 996 44
rect 950 31 952 39
rect 966 35 968 39
rect 959 33 968 35
rect 980 38 986 40
rect 980 36 982 38
rect 984 36 986 38
rect 980 34 986 36
rect 990 39 996 41
rect 990 37 992 39
rect 994 37 996 39
rect 990 35 996 37
rect 959 31 961 33
rect 963 31 968 33
rect 845 19 847 22
rect 817 13 819 18
rect 824 13 826 18
rect 845 17 850 19
rect 848 9 850 17
rect 861 13 863 17
rect 871 9 873 17
rect 909 16 911 20
rect 959 29 968 31
rect 984 31 986 34
rect 966 26 968 29
rect 976 26 978 30
rect 984 29 988 31
rect 986 26 988 29
rect 993 26 995 35
rect 950 19 952 22
rect 881 9 883 14
rect 888 9 890 14
rect 848 7 873 9
rect 922 13 924 18
rect 929 13 931 18
rect 950 17 955 19
rect 953 9 955 17
rect 966 13 968 17
rect 976 9 978 17
rect 986 9 988 14
rect 993 9 995 14
rect 953 7 978 9
<< ndif >>
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 9 22 14 25
rect 16 25 24 31
rect 26 29 34 31
rect 26 27 29 29
rect 31 27 34 29
rect 26 25 34 27
rect 36 25 43 31
rect 88 29 95 31
rect 49 26 54 29
rect 16 22 22 25
rect 18 18 22 22
rect 38 18 43 25
rect 47 24 54 26
rect 47 22 49 24
rect 51 22 54 24
rect 47 20 54 22
rect 56 20 67 29
rect 18 16 24 18
rect 18 14 20 16
rect 22 14 24 16
rect 18 12 24 14
rect 37 16 43 18
rect 58 18 67 20
rect 69 18 74 29
rect 76 24 81 29
rect 88 27 90 29
rect 92 27 95 29
rect 88 25 95 27
rect 76 22 83 24
rect 90 22 95 25
rect 97 26 102 31
rect 193 29 200 31
rect 154 26 159 29
rect 97 22 111 26
rect 76 20 79 22
rect 81 20 83 22
rect 76 18 83 20
rect 102 21 111 22
rect 102 19 104 21
rect 106 19 111 21
rect 37 14 39 16
rect 41 14 43 16
rect 37 12 43 14
rect 58 12 65 18
rect 102 17 111 19
rect 113 24 121 26
rect 113 22 116 24
rect 118 22 121 24
rect 113 17 121 22
rect 123 22 131 26
rect 123 20 126 22
rect 128 20 131 22
rect 123 17 131 20
rect 58 10 60 12
rect 62 10 65 12
rect 58 8 65 10
rect 126 14 131 17
rect 133 14 138 26
rect 140 14 148 26
rect 152 24 159 26
rect 152 22 154 24
rect 156 22 159 24
rect 152 20 159 22
rect 161 20 172 29
rect 163 18 172 20
rect 174 18 179 29
rect 181 24 186 29
rect 193 27 195 29
rect 197 27 200 29
rect 193 25 200 27
rect 181 22 188 24
rect 195 22 200 25
rect 202 26 207 31
rect 257 29 264 31
rect 257 27 259 29
rect 261 27 264 29
rect 202 22 216 26
rect 181 20 184 22
rect 186 20 188 22
rect 181 18 188 20
rect 207 21 216 22
rect 207 19 209 21
rect 211 19 216 21
rect 142 12 148 14
rect 142 10 144 12
rect 146 10 148 12
rect 142 8 148 10
rect 163 12 170 18
rect 207 17 216 19
rect 218 24 226 26
rect 218 22 221 24
rect 223 22 226 24
rect 218 17 226 22
rect 228 22 236 26
rect 228 20 231 22
rect 233 20 236 22
rect 228 17 236 20
rect 163 10 165 12
rect 167 10 170 12
rect 163 8 170 10
rect 231 14 236 17
rect 238 14 243 26
rect 245 14 253 26
rect 257 25 264 27
rect 259 22 264 25
rect 266 25 274 31
rect 276 29 284 31
rect 276 27 279 29
rect 281 27 284 29
rect 276 25 284 27
rect 286 25 293 31
rect 338 29 345 31
rect 299 26 304 29
rect 266 22 272 25
rect 268 18 272 22
rect 288 18 293 25
rect 297 24 304 26
rect 297 22 299 24
rect 301 22 304 24
rect 297 20 304 22
rect 306 20 317 29
rect 268 16 274 18
rect 268 14 270 16
rect 272 14 274 16
rect 247 12 253 14
rect 247 10 249 12
rect 251 10 253 12
rect 247 8 253 10
rect 268 12 274 14
rect 287 16 293 18
rect 308 18 317 20
rect 319 18 324 29
rect 326 24 331 29
rect 338 27 340 29
rect 342 27 345 29
rect 338 25 345 27
rect 326 22 333 24
rect 340 22 345 25
rect 347 26 352 31
rect 443 29 450 31
rect 404 26 409 29
rect 347 22 361 26
rect 326 20 329 22
rect 331 20 333 22
rect 326 18 333 20
rect 352 21 361 22
rect 352 19 354 21
rect 356 19 361 21
rect 287 14 289 16
rect 291 14 293 16
rect 287 12 293 14
rect 308 12 315 18
rect 352 17 361 19
rect 363 24 371 26
rect 363 22 366 24
rect 368 22 371 24
rect 363 17 371 22
rect 373 22 381 26
rect 373 20 376 22
rect 378 20 381 22
rect 373 17 381 20
rect 308 10 310 12
rect 312 10 315 12
rect 308 8 315 10
rect 376 14 381 17
rect 383 14 388 26
rect 390 14 398 26
rect 402 24 409 26
rect 402 22 404 24
rect 406 22 409 24
rect 402 20 409 22
rect 411 20 422 29
rect 413 18 422 20
rect 424 18 429 29
rect 431 24 436 29
rect 443 27 445 29
rect 447 27 450 29
rect 443 25 450 27
rect 431 22 438 24
rect 445 22 450 25
rect 452 26 457 31
rect 507 29 514 31
rect 507 27 509 29
rect 511 27 514 29
rect 452 22 466 26
rect 431 20 434 22
rect 436 20 438 22
rect 431 18 438 20
rect 457 21 466 22
rect 457 19 459 21
rect 461 19 466 21
rect 392 12 398 14
rect 392 10 394 12
rect 396 10 398 12
rect 392 8 398 10
rect 413 12 420 18
rect 457 17 466 19
rect 468 24 476 26
rect 468 22 471 24
rect 473 22 476 24
rect 468 17 476 22
rect 478 22 486 26
rect 478 20 481 22
rect 483 20 486 22
rect 478 17 486 20
rect 413 10 415 12
rect 417 10 420 12
rect 413 8 420 10
rect 481 14 486 17
rect 488 14 493 26
rect 495 14 503 26
rect 507 25 514 27
rect 509 22 514 25
rect 516 25 524 31
rect 526 29 534 31
rect 526 27 529 29
rect 531 27 534 29
rect 526 25 534 27
rect 536 25 543 31
rect 588 29 595 31
rect 549 26 554 29
rect 516 22 522 25
rect 518 18 522 22
rect 538 18 543 25
rect 547 24 554 26
rect 547 22 549 24
rect 551 22 554 24
rect 547 20 554 22
rect 556 20 567 29
rect 518 16 524 18
rect 518 14 520 16
rect 522 14 524 16
rect 497 12 503 14
rect 497 10 499 12
rect 501 10 503 12
rect 497 8 503 10
rect 518 12 524 14
rect 537 16 543 18
rect 558 18 567 20
rect 569 18 574 29
rect 576 24 581 29
rect 588 27 590 29
rect 592 27 595 29
rect 588 25 595 27
rect 576 22 583 24
rect 590 22 595 25
rect 597 26 602 31
rect 693 29 700 31
rect 654 26 659 29
rect 597 22 611 26
rect 576 20 579 22
rect 581 20 583 22
rect 576 18 583 20
rect 602 21 611 22
rect 602 19 604 21
rect 606 19 611 21
rect 537 14 539 16
rect 541 14 543 16
rect 537 12 543 14
rect 558 12 565 18
rect 602 17 611 19
rect 613 24 621 26
rect 613 22 616 24
rect 618 22 621 24
rect 613 17 621 22
rect 623 22 631 26
rect 623 20 626 22
rect 628 20 631 22
rect 623 17 631 20
rect 558 10 560 12
rect 562 10 565 12
rect 558 8 565 10
rect 626 14 631 17
rect 633 14 638 26
rect 640 14 648 26
rect 652 24 659 26
rect 652 22 654 24
rect 656 22 659 24
rect 652 20 659 22
rect 661 20 672 29
rect 663 18 672 20
rect 674 18 679 29
rect 681 24 686 29
rect 693 27 695 29
rect 697 27 700 29
rect 693 25 700 27
rect 681 22 688 24
rect 695 22 700 25
rect 702 26 707 31
rect 757 29 764 31
rect 757 27 759 29
rect 761 27 764 29
rect 702 22 716 26
rect 681 20 684 22
rect 686 20 688 22
rect 681 18 688 20
rect 707 21 716 22
rect 707 19 709 21
rect 711 19 716 21
rect 642 12 648 14
rect 642 10 644 12
rect 646 10 648 12
rect 642 8 648 10
rect 663 12 670 18
rect 707 17 716 19
rect 718 24 726 26
rect 718 22 721 24
rect 723 22 726 24
rect 718 17 726 22
rect 728 22 736 26
rect 728 20 731 22
rect 733 20 736 22
rect 728 17 736 20
rect 663 10 665 12
rect 667 10 670 12
rect 663 8 670 10
rect 731 14 736 17
rect 738 14 743 26
rect 745 14 753 26
rect 757 25 764 27
rect 759 22 764 25
rect 766 25 774 31
rect 776 29 784 31
rect 776 27 779 29
rect 781 27 784 29
rect 776 25 784 27
rect 786 25 793 31
rect 838 29 845 31
rect 799 26 804 29
rect 766 22 772 25
rect 768 18 772 22
rect 788 18 793 25
rect 797 24 804 26
rect 797 22 799 24
rect 801 22 804 24
rect 797 20 804 22
rect 806 20 817 29
rect 768 16 774 18
rect 768 14 770 16
rect 772 14 774 16
rect 747 12 753 14
rect 747 10 749 12
rect 751 10 753 12
rect 747 8 753 10
rect 768 12 774 14
rect 787 16 793 18
rect 808 18 817 20
rect 819 18 824 29
rect 826 24 831 29
rect 838 27 840 29
rect 842 27 845 29
rect 838 25 845 27
rect 826 22 833 24
rect 840 22 845 25
rect 847 26 852 31
rect 943 29 950 31
rect 904 26 909 29
rect 847 22 861 26
rect 826 20 829 22
rect 831 20 833 22
rect 826 18 833 20
rect 852 21 861 22
rect 852 19 854 21
rect 856 19 861 21
rect 787 14 789 16
rect 791 14 793 16
rect 787 12 793 14
rect 808 12 815 18
rect 852 17 861 19
rect 863 24 871 26
rect 863 22 866 24
rect 868 22 871 24
rect 863 17 871 22
rect 873 22 881 26
rect 873 20 876 22
rect 878 20 881 22
rect 873 17 881 20
rect 808 10 810 12
rect 812 10 815 12
rect 808 8 815 10
rect 876 14 881 17
rect 883 14 888 26
rect 890 14 898 26
rect 902 24 909 26
rect 902 22 904 24
rect 906 22 909 24
rect 902 20 909 22
rect 911 20 922 29
rect 913 18 922 20
rect 924 18 929 29
rect 931 24 936 29
rect 943 27 945 29
rect 947 27 950 29
rect 943 25 950 27
rect 931 22 938 24
rect 945 22 950 25
rect 952 26 957 31
rect 952 22 966 26
rect 931 20 934 22
rect 936 20 938 22
rect 931 18 938 20
rect 957 21 966 22
rect 957 19 959 21
rect 961 19 966 21
rect 892 12 898 14
rect 892 10 894 12
rect 896 10 898 12
rect 892 8 898 10
rect 913 12 920 18
rect 957 17 966 19
rect 968 24 976 26
rect 968 22 971 24
rect 973 22 976 24
rect 968 17 976 22
rect 978 22 986 26
rect 978 20 981 22
rect 983 20 986 22
rect 978 17 986 20
rect 913 10 915 12
rect 917 10 920 12
rect 913 8 920 10
rect 981 14 986 17
rect 988 14 993 26
rect 995 14 1003 26
rect 997 12 1003 14
rect 997 10 999 12
rect 1001 10 1003 12
rect 997 8 1003 10
<< pdif >>
rect 18 69 27 71
rect 18 67 20 69
rect 22 67 27 69
rect 18 61 27 67
rect 7 59 14 61
rect 7 57 9 59
rect 11 57 14 59
rect 7 52 14 57
rect 7 50 9 52
rect 11 50 14 52
rect 7 48 14 50
rect 9 43 14 48
rect 16 50 27 61
rect 29 50 34 71
rect 36 64 41 71
rect 36 62 43 64
rect 58 62 64 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 58 43 60
rect 36 50 41 58
rect 49 57 54 62
rect 47 55 54 57
rect 47 53 49 55
rect 51 53 54 55
rect 16 43 24 50
rect 47 48 54 53
rect 47 46 49 48
rect 51 46 54 48
rect 47 44 54 46
rect 56 60 64 62
rect 56 58 59 60
rect 61 58 64 60
rect 56 51 64 58
rect 66 62 74 64
rect 66 60 69 62
rect 71 60 74 62
rect 66 55 74 60
rect 66 53 69 55
rect 71 53 74 55
rect 66 51 74 53
rect 76 62 83 64
rect 76 60 79 62
rect 81 60 83 62
rect 76 51 83 60
rect 56 44 62 51
rect 98 50 103 71
rect 96 48 103 50
rect 96 46 98 48
rect 100 46 103 48
rect 96 44 103 46
rect 105 69 117 71
rect 105 67 108 69
rect 110 67 117 69
rect 105 62 117 67
rect 134 62 139 71
rect 105 60 108 62
rect 110 60 119 62
rect 105 44 119 60
rect 121 55 129 62
rect 121 53 124 55
rect 126 53 129 55
rect 121 48 129 53
rect 121 46 124 48
rect 126 46 129 48
rect 121 44 129 46
rect 131 55 139 62
rect 131 53 134 55
rect 136 53 139 55
rect 131 44 139 53
rect 141 65 146 71
rect 141 63 148 65
rect 141 61 144 63
rect 146 61 148 63
rect 163 62 169 64
rect 141 59 148 61
rect 141 44 146 59
rect 154 57 159 62
rect 152 55 159 57
rect 152 53 154 55
rect 156 53 159 55
rect 152 48 159 53
rect 152 46 154 48
rect 156 46 159 48
rect 152 44 159 46
rect 161 60 169 62
rect 161 58 164 60
rect 166 58 169 60
rect 161 51 169 58
rect 171 62 179 64
rect 171 60 174 62
rect 176 60 179 62
rect 171 55 179 60
rect 171 53 174 55
rect 176 53 179 55
rect 171 51 179 53
rect 181 62 188 64
rect 181 60 184 62
rect 186 60 188 62
rect 181 51 188 60
rect 161 44 167 51
rect 203 50 208 71
rect 201 48 208 50
rect 201 46 203 48
rect 205 46 208 48
rect 201 44 208 46
rect 210 69 222 71
rect 210 67 213 69
rect 215 67 222 69
rect 210 62 222 67
rect 239 62 244 71
rect 210 60 213 62
rect 215 60 224 62
rect 210 44 224 60
rect 226 55 234 62
rect 226 53 229 55
rect 231 53 234 55
rect 226 48 234 53
rect 226 46 229 48
rect 231 46 234 48
rect 226 44 234 46
rect 236 55 244 62
rect 236 53 239 55
rect 241 53 244 55
rect 236 44 244 53
rect 246 65 251 71
rect 268 69 277 71
rect 268 67 270 69
rect 272 67 277 69
rect 246 63 253 65
rect 246 61 249 63
rect 251 61 253 63
rect 268 61 277 67
rect 246 59 253 61
rect 257 59 264 61
rect 246 44 251 59
rect 257 57 259 59
rect 261 57 264 59
rect 257 52 264 57
rect 257 50 259 52
rect 261 50 264 52
rect 257 48 264 50
rect 259 43 264 48
rect 266 50 277 61
rect 279 50 284 71
rect 286 64 291 71
rect 286 62 293 64
rect 308 62 314 64
rect 286 60 289 62
rect 291 60 293 62
rect 286 58 293 60
rect 286 50 291 58
rect 299 57 304 62
rect 297 55 304 57
rect 297 53 299 55
rect 301 53 304 55
rect 266 43 274 50
rect 297 48 304 53
rect 297 46 299 48
rect 301 46 304 48
rect 297 44 304 46
rect 306 60 314 62
rect 306 58 309 60
rect 311 58 314 60
rect 306 51 314 58
rect 316 62 324 64
rect 316 60 319 62
rect 321 60 324 62
rect 316 55 324 60
rect 316 53 319 55
rect 321 53 324 55
rect 316 51 324 53
rect 326 62 333 64
rect 326 60 329 62
rect 331 60 333 62
rect 326 51 333 60
rect 306 44 312 51
rect 348 50 353 71
rect 346 48 353 50
rect 346 46 348 48
rect 350 46 353 48
rect 346 44 353 46
rect 355 69 367 71
rect 355 67 358 69
rect 360 67 367 69
rect 355 62 367 67
rect 384 62 389 71
rect 355 60 358 62
rect 360 60 369 62
rect 355 44 369 60
rect 371 55 379 62
rect 371 53 374 55
rect 376 53 379 55
rect 371 48 379 53
rect 371 46 374 48
rect 376 46 379 48
rect 371 44 379 46
rect 381 55 389 62
rect 381 53 384 55
rect 386 53 389 55
rect 381 44 389 53
rect 391 65 396 71
rect 391 63 398 65
rect 391 61 394 63
rect 396 61 398 63
rect 413 62 419 64
rect 391 59 398 61
rect 391 44 396 59
rect 404 57 409 62
rect 402 55 409 57
rect 402 53 404 55
rect 406 53 409 55
rect 402 48 409 53
rect 402 46 404 48
rect 406 46 409 48
rect 402 44 409 46
rect 411 60 419 62
rect 411 58 414 60
rect 416 58 419 60
rect 411 51 419 58
rect 421 62 429 64
rect 421 60 424 62
rect 426 60 429 62
rect 421 55 429 60
rect 421 53 424 55
rect 426 53 429 55
rect 421 51 429 53
rect 431 62 438 64
rect 431 60 434 62
rect 436 60 438 62
rect 431 51 438 60
rect 411 44 417 51
rect 453 50 458 71
rect 451 48 458 50
rect 451 46 453 48
rect 455 46 458 48
rect 451 44 458 46
rect 460 69 472 71
rect 460 67 463 69
rect 465 67 472 69
rect 460 62 472 67
rect 489 62 494 71
rect 460 60 463 62
rect 465 60 474 62
rect 460 44 474 60
rect 476 55 484 62
rect 476 53 479 55
rect 481 53 484 55
rect 476 48 484 53
rect 476 46 479 48
rect 481 46 484 48
rect 476 44 484 46
rect 486 55 494 62
rect 486 53 489 55
rect 491 53 494 55
rect 486 44 494 53
rect 496 65 501 71
rect 518 69 527 71
rect 518 67 520 69
rect 522 67 527 69
rect 496 63 503 65
rect 496 61 499 63
rect 501 61 503 63
rect 518 61 527 67
rect 496 59 503 61
rect 507 59 514 61
rect 496 44 501 59
rect 507 57 509 59
rect 511 57 514 59
rect 507 52 514 57
rect 507 50 509 52
rect 511 50 514 52
rect 507 48 514 50
rect 509 43 514 48
rect 516 50 527 61
rect 529 50 534 71
rect 536 64 541 71
rect 536 62 543 64
rect 558 62 564 64
rect 536 60 539 62
rect 541 60 543 62
rect 536 58 543 60
rect 536 50 541 58
rect 549 57 554 62
rect 547 55 554 57
rect 547 53 549 55
rect 551 53 554 55
rect 516 43 524 50
rect 547 48 554 53
rect 547 46 549 48
rect 551 46 554 48
rect 547 44 554 46
rect 556 60 564 62
rect 556 58 559 60
rect 561 58 564 60
rect 556 51 564 58
rect 566 62 574 64
rect 566 60 569 62
rect 571 60 574 62
rect 566 55 574 60
rect 566 53 569 55
rect 571 53 574 55
rect 566 51 574 53
rect 576 62 583 64
rect 576 60 579 62
rect 581 60 583 62
rect 576 51 583 60
rect 556 44 562 51
rect 598 50 603 71
rect 596 48 603 50
rect 596 46 598 48
rect 600 46 603 48
rect 596 44 603 46
rect 605 69 617 71
rect 605 67 608 69
rect 610 67 617 69
rect 605 62 617 67
rect 634 62 639 71
rect 605 60 608 62
rect 610 60 619 62
rect 605 44 619 60
rect 621 55 629 62
rect 621 53 624 55
rect 626 53 629 55
rect 621 48 629 53
rect 621 46 624 48
rect 626 46 629 48
rect 621 44 629 46
rect 631 55 639 62
rect 631 53 634 55
rect 636 53 639 55
rect 631 44 639 53
rect 641 65 646 71
rect 641 63 648 65
rect 641 61 644 63
rect 646 61 648 63
rect 663 62 669 64
rect 641 59 648 61
rect 641 44 646 59
rect 654 57 659 62
rect 652 55 659 57
rect 652 53 654 55
rect 656 53 659 55
rect 652 48 659 53
rect 652 46 654 48
rect 656 46 659 48
rect 652 44 659 46
rect 661 60 669 62
rect 661 58 664 60
rect 666 58 669 60
rect 661 51 669 58
rect 671 62 679 64
rect 671 60 674 62
rect 676 60 679 62
rect 671 55 679 60
rect 671 53 674 55
rect 676 53 679 55
rect 671 51 679 53
rect 681 62 688 64
rect 681 60 684 62
rect 686 60 688 62
rect 681 51 688 60
rect 661 44 667 51
rect 703 50 708 71
rect 701 48 708 50
rect 701 46 703 48
rect 705 46 708 48
rect 701 44 708 46
rect 710 69 722 71
rect 710 67 713 69
rect 715 67 722 69
rect 710 62 722 67
rect 739 62 744 71
rect 710 60 713 62
rect 715 60 724 62
rect 710 44 724 60
rect 726 55 734 62
rect 726 53 729 55
rect 731 53 734 55
rect 726 48 734 53
rect 726 46 729 48
rect 731 46 734 48
rect 726 44 734 46
rect 736 55 744 62
rect 736 53 739 55
rect 741 53 744 55
rect 736 44 744 53
rect 746 65 751 71
rect 768 69 777 71
rect 768 67 770 69
rect 772 67 777 69
rect 746 63 753 65
rect 746 61 749 63
rect 751 61 753 63
rect 768 61 777 67
rect 746 59 753 61
rect 757 59 764 61
rect 746 44 751 59
rect 757 57 759 59
rect 761 57 764 59
rect 757 52 764 57
rect 757 50 759 52
rect 761 50 764 52
rect 757 48 764 50
rect 759 43 764 48
rect 766 50 777 61
rect 779 50 784 71
rect 786 64 791 71
rect 786 62 793 64
rect 808 62 814 64
rect 786 60 789 62
rect 791 60 793 62
rect 786 58 793 60
rect 786 50 791 58
rect 799 57 804 62
rect 797 55 804 57
rect 797 53 799 55
rect 801 53 804 55
rect 766 43 774 50
rect 797 48 804 53
rect 797 46 799 48
rect 801 46 804 48
rect 797 44 804 46
rect 806 60 814 62
rect 806 58 809 60
rect 811 58 814 60
rect 806 51 814 58
rect 816 62 824 64
rect 816 60 819 62
rect 821 60 824 62
rect 816 55 824 60
rect 816 53 819 55
rect 821 53 824 55
rect 816 51 824 53
rect 826 62 833 64
rect 826 60 829 62
rect 831 60 833 62
rect 826 51 833 60
rect 806 44 812 51
rect 848 50 853 71
rect 846 48 853 50
rect 846 46 848 48
rect 850 46 853 48
rect 846 44 853 46
rect 855 69 867 71
rect 855 67 858 69
rect 860 67 867 69
rect 855 62 867 67
rect 884 62 889 71
rect 855 60 858 62
rect 860 60 869 62
rect 855 44 869 60
rect 871 55 879 62
rect 871 53 874 55
rect 876 53 879 55
rect 871 48 879 53
rect 871 46 874 48
rect 876 46 879 48
rect 871 44 879 46
rect 881 55 889 62
rect 881 53 884 55
rect 886 53 889 55
rect 881 44 889 53
rect 891 65 896 71
rect 891 63 898 65
rect 891 61 894 63
rect 896 61 898 63
rect 913 62 919 64
rect 891 59 898 61
rect 891 44 896 59
rect 904 57 909 62
rect 902 55 909 57
rect 902 53 904 55
rect 906 53 909 55
rect 902 48 909 53
rect 902 46 904 48
rect 906 46 909 48
rect 902 44 909 46
rect 911 60 919 62
rect 911 58 914 60
rect 916 58 919 60
rect 911 51 919 58
rect 921 62 929 64
rect 921 60 924 62
rect 926 60 929 62
rect 921 55 929 60
rect 921 53 924 55
rect 926 53 929 55
rect 921 51 929 53
rect 931 62 938 64
rect 931 60 934 62
rect 936 60 938 62
rect 931 51 938 60
rect 911 44 917 51
rect 953 50 958 71
rect 951 48 958 50
rect 951 46 953 48
rect 955 46 958 48
rect 951 44 958 46
rect 960 69 972 71
rect 960 67 963 69
rect 965 67 972 69
rect 960 62 972 67
rect 989 62 994 71
rect 960 60 963 62
rect 965 60 974 62
rect 960 44 974 60
rect 976 55 984 62
rect 976 53 979 55
rect 981 53 984 55
rect 976 48 984 53
rect 976 46 979 48
rect 981 46 984 48
rect 976 44 984 46
rect 986 55 994 62
rect 986 53 989 55
rect 991 53 994 55
rect 986 44 994 53
rect 996 65 1001 71
rect 996 63 1003 65
rect 996 61 999 63
rect 1001 61 1003 63
rect 996 59 1003 61
rect 996 44 1001 59
<< alu1 >>
rect 3 72 1007 77
rect 3 70 10 72
rect 12 70 50 72
rect 52 70 124 72
rect 126 70 155 72
rect 157 70 229 72
rect 231 70 260 72
rect 262 70 300 72
rect 302 70 374 72
rect 376 70 405 72
rect 407 70 479 72
rect 481 70 510 72
rect 512 70 550 72
rect 552 70 624 72
rect 626 70 655 72
rect 657 70 729 72
rect 731 70 760 72
rect 762 70 800 72
rect 802 70 874 72
rect 876 70 905 72
rect 907 70 979 72
rect 981 70 1007 72
rect 3 69 1007 70
rect 7 63 11 64
rect 7 59 20 63
rect 7 57 9 59
rect 7 52 11 57
rect 7 50 9 52
rect 7 31 11 50
rect 39 55 43 56
rect 39 53 40 55
rect 42 53 43 55
rect 39 47 43 53
rect 22 45 43 47
rect 22 43 36 45
rect 38 43 43 45
rect 47 55 52 57
rect 47 53 49 55
rect 51 53 52 55
rect 88 58 100 64
rect 47 48 52 53
rect 47 46 49 48
rect 51 46 52 48
rect 47 44 52 46
rect 47 39 51 44
rect 7 29 12 31
rect 7 27 9 29
rect 11 27 12 29
rect 7 25 12 27
rect 22 38 51 39
rect 22 36 26 38
rect 28 36 51 38
rect 22 35 51 36
rect 39 26 43 35
rect 47 24 51 35
rect 79 49 83 56
rect 88 49 93 58
rect 79 47 93 49
rect 70 46 93 47
rect 70 44 76 46
rect 78 44 90 46
rect 92 44 93 46
rect 70 43 83 44
rect 87 43 93 44
rect 88 42 93 43
rect 62 38 76 39
rect 62 36 66 38
rect 68 36 76 38
rect 62 35 76 36
rect 47 22 49 24
rect 51 22 59 24
rect 47 18 59 22
rect 71 29 76 35
rect 71 27 72 29
rect 74 27 76 29
rect 71 26 76 27
rect 104 33 109 40
rect 132 55 148 56
rect 132 53 134 55
rect 136 53 148 55
rect 132 51 148 53
rect 104 32 106 33
rect 96 31 106 32
rect 108 31 109 33
rect 96 29 109 31
rect 96 27 99 29
rect 101 27 109 29
rect 96 26 109 27
rect 144 29 148 51
rect 144 27 145 29
rect 147 27 148 29
rect 144 23 148 27
rect 124 22 148 23
rect 124 20 126 22
rect 128 20 148 22
rect 124 19 148 20
rect 152 55 157 57
rect 152 53 154 55
rect 156 53 157 55
rect 193 58 205 64
rect 257 63 261 64
rect 152 48 157 53
rect 152 46 154 48
rect 156 46 157 48
rect 152 44 157 46
rect 152 24 156 44
rect 184 49 188 56
rect 193 49 198 58
rect 257 59 270 63
rect 257 57 259 59
rect 184 47 198 49
rect 175 46 187 47
rect 175 44 181 46
rect 183 45 187 46
rect 189 46 198 47
rect 189 45 195 46
rect 183 44 195 45
rect 197 44 198 46
rect 175 43 188 44
rect 192 43 198 44
rect 193 42 198 43
rect 167 38 181 39
rect 167 36 171 38
rect 173 36 181 38
rect 167 35 181 36
rect 152 22 154 24
rect 156 22 164 24
rect 152 18 164 22
rect 176 29 181 35
rect 176 27 177 29
rect 179 27 181 29
rect 176 26 181 27
rect 209 33 214 40
rect 237 55 253 56
rect 237 53 239 55
rect 241 53 253 55
rect 237 51 253 53
rect 209 32 211 33
rect 201 31 211 32
rect 213 31 214 33
rect 201 29 214 31
rect 201 27 204 29
rect 206 27 214 29
rect 201 26 214 27
rect 249 23 253 51
rect 257 52 261 57
rect 257 50 259 52
rect 257 47 261 50
rect 289 55 293 56
rect 289 53 290 55
rect 292 53 293 55
rect 257 45 258 47
rect 260 45 261 47
rect 257 31 261 45
rect 289 47 293 53
rect 272 45 293 47
rect 272 43 286 45
rect 288 43 293 45
rect 297 55 302 57
rect 297 53 299 55
rect 301 53 302 55
rect 338 58 350 64
rect 297 48 302 53
rect 297 46 299 48
rect 301 46 302 48
rect 297 44 302 46
rect 297 39 301 44
rect 257 29 262 31
rect 257 27 259 29
rect 261 27 262 29
rect 257 25 262 27
rect 272 38 301 39
rect 272 36 276 38
rect 278 36 301 38
rect 272 35 301 36
rect 289 26 293 35
rect 229 22 253 23
rect 229 20 231 22
rect 233 20 253 22
rect 229 19 253 20
rect 297 24 301 35
rect 329 49 333 56
rect 338 49 343 58
rect 329 47 343 49
rect 320 46 343 47
rect 320 44 326 46
rect 328 44 340 46
rect 342 44 343 46
rect 320 43 333 44
rect 337 43 343 44
rect 338 42 343 43
rect 312 38 326 39
rect 312 36 316 38
rect 318 36 326 38
rect 312 35 326 36
rect 297 22 299 24
rect 301 22 309 24
rect 297 18 309 22
rect 321 29 326 35
rect 321 27 322 29
rect 324 27 326 29
rect 321 26 326 27
rect 354 33 359 40
rect 382 55 398 56
rect 382 53 384 55
rect 386 53 398 55
rect 382 51 398 53
rect 354 32 356 33
rect 346 31 356 32
rect 358 31 359 33
rect 346 29 359 31
rect 346 27 349 29
rect 351 27 359 29
rect 346 26 359 27
rect 394 29 398 51
rect 394 27 395 29
rect 397 27 398 29
rect 394 23 398 27
rect 374 22 398 23
rect 374 20 376 22
rect 378 20 398 22
rect 374 19 398 20
rect 402 55 407 57
rect 402 53 404 55
rect 406 53 407 55
rect 443 58 455 64
rect 507 63 511 64
rect 402 48 407 53
rect 402 46 404 48
rect 406 46 407 48
rect 402 44 407 46
rect 402 24 406 44
rect 434 49 438 56
rect 443 49 448 58
rect 507 59 520 63
rect 507 57 509 59
rect 434 47 448 49
rect 425 46 439 47
rect 425 44 431 46
rect 433 45 439 46
rect 441 46 448 47
rect 441 45 445 46
rect 433 44 445 45
rect 447 44 448 46
rect 425 43 438 44
rect 442 43 448 44
rect 443 42 448 43
rect 417 38 431 39
rect 417 36 421 38
rect 423 36 431 38
rect 417 35 431 36
rect 402 22 404 24
rect 406 22 414 24
rect 402 18 414 22
rect 426 29 431 35
rect 426 27 427 29
rect 429 27 431 29
rect 426 26 431 27
rect 459 33 464 40
rect 487 55 503 56
rect 487 53 489 55
rect 491 53 503 55
rect 487 51 503 53
rect 459 32 461 33
rect 451 31 461 32
rect 463 31 464 33
rect 451 29 464 31
rect 451 27 454 29
rect 456 27 464 29
rect 451 26 464 27
rect 499 23 503 51
rect 507 52 511 57
rect 507 50 509 52
rect 507 47 511 50
rect 539 55 543 56
rect 539 53 540 55
rect 542 53 543 55
rect 507 45 508 47
rect 510 45 511 47
rect 507 31 511 45
rect 539 47 543 53
rect 522 45 543 47
rect 522 43 536 45
rect 538 43 543 45
rect 547 55 552 57
rect 547 53 549 55
rect 551 53 552 55
rect 588 58 600 64
rect 547 48 552 53
rect 547 46 549 48
rect 551 46 552 48
rect 547 44 552 46
rect 547 39 551 44
rect 507 29 512 31
rect 507 27 509 29
rect 511 27 512 29
rect 507 25 512 27
rect 522 38 551 39
rect 522 36 526 38
rect 528 36 551 38
rect 522 35 551 36
rect 539 26 543 35
rect 479 22 503 23
rect 479 20 481 22
rect 483 20 503 22
rect 479 19 503 20
rect 547 24 551 35
rect 579 49 583 56
rect 588 49 593 58
rect 579 47 593 49
rect 570 46 593 47
rect 570 44 576 46
rect 578 44 590 46
rect 592 44 593 46
rect 570 43 583 44
rect 587 43 593 44
rect 588 42 593 43
rect 562 38 576 39
rect 562 36 566 38
rect 568 36 576 38
rect 562 35 576 36
rect 547 22 549 24
rect 551 22 559 24
rect 547 18 559 22
rect 571 29 576 35
rect 571 27 572 29
rect 574 27 576 29
rect 571 26 576 27
rect 604 33 609 40
rect 632 55 648 56
rect 632 53 634 55
rect 636 53 648 55
rect 632 51 648 53
rect 604 32 606 33
rect 596 31 606 32
rect 608 31 609 33
rect 596 29 609 31
rect 596 27 599 29
rect 601 27 609 29
rect 596 26 609 27
rect 644 29 648 51
rect 644 27 645 29
rect 647 27 648 29
rect 644 23 648 27
rect 624 22 648 23
rect 624 20 626 22
rect 628 20 648 22
rect 624 19 648 20
rect 652 55 657 57
rect 652 53 654 55
rect 656 53 657 55
rect 693 58 705 64
rect 757 63 761 64
rect 652 48 657 53
rect 652 46 654 48
rect 656 46 657 48
rect 652 44 657 46
rect 652 24 656 44
rect 684 49 688 56
rect 693 49 698 58
rect 757 59 770 63
rect 757 57 759 59
rect 684 47 698 49
rect 675 46 689 47
rect 675 44 681 46
rect 683 45 689 46
rect 691 46 698 47
rect 691 45 695 46
rect 683 44 695 45
rect 697 44 698 46
rect 675 43 688 44
rect 692 43 698 44
rect 693 42 698 43
rect 667 38 681 39
rect 667 36 671 38
rect 673 36 681 38
rect 667 35 681 36
rect 652 22 654 24
rect 656 22 664 24
rect 652 18 664 22
rect 676 29 681 35
rect 676 27 677 29
rect 679 27 681 29
rect 676 26 681 27
rect 709 33 714 40
rect 737 55 753 56
rect 737 53 739 55
rect 741 53 753 55
rect 737 51 753 53
rect 709 32 711 33
rect 701 31 711 32
rect 713 31 714 33
rect 701 29 714 31
rect 701 27 704 29
rect 706 27 714 29
rect 701 26 714 27
rect 749 23 753 51
rect 757 52 761 57
rect 757 50 759 52
rect 757 47 761 50
rect 789 55 793 56
rect 789 53 790 55
rect 792 53 793 55
rect 757 45 758 47
rect 760 45 761 47
rect 757 31 761 45
rect 789 47 793 53
rect 772 45 793 47
rect 772 43 786 45
rect 788 43 793 45
rect 797 55 802 57
rect 797 53 799 55
rect 801 53 802 55
rect 838 58 850 64
rect 797 48 802 53
rect 797 46 799 48
rect 801 46 802 48
rect 797 44 802 46
rect 797 39 801 44
rect 757 29 762 31
rect 757 27 759 29
rect 761 27 762 29
rect 757 25 762 27
rect 772 38 801 39
rect 772 36 776 38
rect 778 36 801 38
rect 772 35 801 36
rect 789 26 793 35
rect 729 22 753 23
rect 729 20 731 22
rect 733 20 753 22
rect 729 19 753 20
rect 797 24 801 35
rect 829 49 833 56
rect 838 49 843 58
rect 829 47 843 49
rect 820 46 843 47
rect 820 44 826 46
rect 828 44 840 46
rect 842 44 843 46
rect 820 43 833 44
rect 837 43 843 44
rect 838 42 843 43
rect 812 38 826 39
rect 812 36 816 38
rect 818 36 826 38
rect 812 35 826 36
rect 797 22 799 24
rect 801 22 809 24
rect 797 18 809 22
rect 821 29 826 35
rect 821 27 822 29
rect 824 27 826 29
rect 821 26 826 27
rect 854 33 859 40
rect 882 55 898 56
rect 882 53 884 55
rect 886 53 898 55
rect 882 51 898 53
rect 854 32 856 33
rect 846 31 856 32
rect 858 31 859 33
rect 846 29 859 31
rect 846 27 849 29
rect 851 27 859 29
rect 846 26 859 27
rect 894 29 898 51
rect 894 27 895 29
rect 897 27 898 29
rect 894 23 898 27
rect 874 22 898 23
rect 874 20 876 22
rect 878 20 898 22
rect 874 19 898 20
rect 902 55 907 57
rect 902 53 904 55
rect 906 53 907 55
rect 943 58 955 64
rect 902 48 907 53
rect 902 46 904 48
rect 906 46 907 48
rect 902 44 907 46
rect 902 24 906 44
rect 934 49 938 56
rect 943 49 948 58
rect 934 47 948 49
rect 925 46 948 47
rect 925 44 931 46
rect 933 44 939 46
rect 941 44 945 46
rect 947 44 948 46
rect 925 43 948 44
rect 943 42 948 43
rect 917 38 931 39
rect 917 36 921 38
rect 923 36 931 38
rect 917 35 931 36
rect 902 22 904 24
rect 906 22 914 24
rect 902 18 914 22
rect 926 29 931 35
rect 926 27 927 29
rect 929 27 931 29
rect 926 26 931 27
rect 959 33 964 40
rect 987 55 1003 56
rect 987 53 989 55
rect 991 53 1003 55
rect 987 51 1003 53
rect 959 32 961 33
rect 951 31 961 32
rect 963 31 964 33
rect 951 29 964 31
rect 951 27 954 29
rect 956 27 964 29
rect 951 26 964 27
rect 999 23 1003 51
rect 979 22 1003 23
rect 979 20 981 22
rect 983 20 1003 22
rect 979 19 1003 20
rect 3 12 1007 13
rect 3 10 10 12
rect 12 10 50 12
rect 52 10 60 12
rect 62 10 91 12
rect 93 10 144 12
rect 146 10 155 12
rect 157 10 165 12
rect 167 10 196 12
rect 198 10 249 12
rect 251 10 260 12
rect 262 10 300 12
rect 302 10 310 12
rect 312 10 341 12
rect 343 10 394 12
rect 396 10 405 12
rect 407 10 415 12
rect 417 10 446 12
rect 448 10 499 12
rect 501 10 510 12
rect 512 10 550 12
rect 552 10 560 12
rect 562 10 591 12
rect 593 10 644 12
rect 646 10 655 12
rect 657 10 665 12
rect 667 10 696 12
rect 698 10 749 12
rect 751 10 760 12
rect 762 10 800 12
rect 802 10 810 12
rect 812 10 841 12
rect 843 10 894 12
rect 896 10 905 12
rect 907 10 915 12
rect 917 11 946 12
rect 917 10 939 11
rect 3 9 939 10
rect 941 10 946 11
rect 948 10 999 12
rect 1001 10 1007 12
rect 941 9 1007 10
rect 3 5 1007 9
<< alu2 >>
rect 39 55 157 56
rect 39 53 40 55
rect 42 53 154 55
rect 156 53 157 55
rect 39 52 157 53
rect 289 55 407 56
rect 289 53 290 55
rect 292 53 404 55
rect 406 53 407 55
rect 289 52 407 53
rect 539 55 657 56
rect 539 53 540 55
rect 542 53 654 55
rect 656 53 657 55
rect 539 52 657 53
rect 789 55 907 56
rect 789 53 790 55
rect 792 53 904 55
rect 906 53 907 55
rect 789 52 907 53
rect 186 47 261 48
rect 186 45 187 47
rect 189 45 258 47
rect 260 45 261 47
rect 186 44 261 45
rect 438 47 511 48
rect 438 45 439 47
rect 441 45 508 47
rect 510 45 511 47
rect 438 44 511 45
rect 688 47 761 48
rect 688 45 689 47
rect 691 45 758 47
rect 760 45 761 47
rect 688 44 761 45
rect 938 46 942 47
rect 938 44 939 46
rect 941 44 942 46
rect 938 37 942 44
rect 938 35 939 37
rect 941 35 942 37
rect 938 34 942 35
rect 71 29 104 30
rect 71 27 72 29
rect 74 27 99 29
rect 101 27 104 29
rect 71 26 104 27
rect 144 29 209 30
rect 144 27 145 29
rect 147 27 177 29
rect 179 27 204 29
rect 206 27 209 29
rect 144 26 209 27
rect 321 29 354 30
rect 321 27 322 29
rect 324 27 349 29
rect 351 27 354 29
rect 321 26 354 27
rect 394 29 459 30
rect 394 27 395 29
rect 397 27 427 29
rect 429 27 454 29
rect 456 27 459 29
rect 394 26 459 27
rect 571 29 604 30
rect 571 27 572 29
rect 574 27 599 29
rect 601 27 604 29
rect 571 26 604 27
rect 644 29 709 30
rect 644 27 645 29
rect 647 27 677 29
rect 679 27 704 29
rect 706 27 709 29
rect 644 26 709 27
rect 821 29 854 30
rect 821 27 822 29
rect 824 27 849 29
rect 851 27 854 29
rect 821 26 854 27
rect 894 29 959 30
rect 894 27 895 29
rect 897 27 927 29
rect 929 27 954 29
rect 956 27 959 29
rect 894 26 959 27
rect 938 21 942 22
rect 938 19 939 21
rect 941 19 942 21
rect 938 11 942 19
rect 938 9 939 11
rect 941 9 942 11
rect 938 7 942 9
<< alu3 >>
rect 938 37 942 38
rect 938 35 939 37
rect 941 35 942 37
rect 938 21 942 35
rect 938 19 939 21
rect 941 19 942 21
rect 938 18 942 19
<< ptie >>
rect 8 12 14 14
rect 48 12 54 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 48 10 50 12
rect 52 10 54 12
rect 48 8 54 10
rect 89 12 95 14
rect 89 10 91 12
rect 93 10 95 12
rect 89 8 95 10
rect 153 12 159 14
rect 153 10 155 12
rect 157 10 159 12
rect 153 8 159 10
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
rect 258 12 264 14
rect 298 12 304 14
rect 258 10 260 12
rect 262 10 264 12
rect 258 8 264 10
rect 298 10 300 12
rect 302 10 304 12
rect 298 8 304 10
rect 339 12 345 14
rect 339 10 341 12
rect 343 10 345 12
rect 339 8 345 10
rect 403 12 409 14
rect 403 10 405 12
rect 407 10 409 12
rect 403 8 409 10
rect 444 12 450 14
rect 444 10 446 12
rect 448 10 450 12
rect 444 8 450 10
rect 508 12 514 14
rect 548 12 554 14
rect 508 10 510 12
rect 512 10 514 12
rect 508 8 514 10
rect 548 10 550 12
rect 552 10 554 12
rect 548 8 554 10
rect 589 12 595 14
rect 589 10 591 12
rect 593 10 595 12
rect 589 8 595 10
rect 653 12 659 14
rect 653 10 655 12
rect 657 10 659 12
rect 653 8 659 10
rect 694 12 700 14
rect 694 10 696 12
rect 698 10 700 12
rect 694 8 700 10
rect 758 12 764 14
rect 798 12 804 14
rect 758 10 760 12
rect 762 10 764 12
rect 758 8 764 10
rect 798 10 800 12
rect 802 10 804 12
rect 798 8 804 10
rect 839 12 845 14
rect 839 10 841 12
rect 843 10 845 12
rect 839 8 845 10
rect 903 12 909 14
rect 903 10 905 12
rect 907 10 909 12
rect 903 8 909 10
rect 944 12 950 14
rect 944 10 946 12
rect 948 10 950 12
rect 944 8 950 10
<< ntie >>
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 48 72 54 74
rect 8 68 14 70
rect 48 70 50 72
rect 52 70 54 72
rect 122 72 128 74
rect 48 68 54 70
rect 122 70 124 72
rect 126 70 128 72
rect 153 72 159 74
rect 122 68 128 70
rect 153 70 155 72
rect 157 70 159 72
rect 227 72 233 74
rect 153 68 159 70
rect 227 70 229 72
rect 231 70 233 72
rect 258 72 264 74
rect 227 68 233 70
rect 258 70 260 72
rect 262 70 264 72
rect 298 72 304 74
rect 258 68 264 70
rect 298 70 300 72
rect 302 70 304 72
rect 372 72 378 74
rect 298 68 304 70
rect 372 70 374 72
rect 376 70 378 72
rect 403 72 409 74
rect 372 68 378 70
rect 403 70 405 72
rect 407 70 409 72
rect 477 72 483 74
rect 403 68 409 70
rect 477 70 479 72
rect 481 70 483 72
rect 508 72 514 74
rect 477 68 483 70
rect 508 70 510 72
rect 512 70 514 72
rect 548 72 554 74
rect 508 68 514 70
rect 548 70 550 72
rect 552 70 554 72
rect 622 72 628 74
rect 548 68 554 70
rect 622 70 624 72
rect 626 70 628 72
rect 653 72 659 74
rect 622 68 628 70
rect 653 70 655 72
rect 657 70 659 72
rect 727 72 733 74
rect 653 68 659 70
rect 727 70 729 72
rect 731 70 733 72
rect 758 72 764 74
rect 727 68 733 70
rect 758 70 760 72
rect 762 70 764 72
rect 798 72 804 74
rect 758 68 764 70
rect 798 70 800 72
rect 802 70 804 72
rect 872 72 878 74
rect 798 68 804 70
rect 872 70 874 72
rect 876 70 878 72
rect 903 72 909 74
rect 872 68 878 70
rect 903 70 905 72
rect 907 70 909 72
rect 977 72 983 74
rect 903 68 909 70
rect 977 70 979 72
rect 981 70 983 72
rect 977 68 983 70
<< nmos >>
rect 14 22 16 31
rect 24 25 26 31
rect 34 25 36 31
rect 54 20 56 29
rect 67 18 69 29
rect 74 18 76 29
rect 95 22 97 31
rect 111 17 113 26
rect 121 17 123 26
rect 131 14 133 26
rect 138 14 140 26
rect 159 20 161 29
rect 172 18 174 29
rect 179 18 181 29
rect 200 22 202 31
rect 216 17 218 26
rect 226 17 228 26
rect 236 14 238 26
rect 243 14 245 26
rect 264 22 266 31
rect 274 25 276 31
rect 284 25 286 31
rect 304 20 306 29
rect 317 18 319 29
rect 324 18 326 29
rect 345 22 347 31
rect 361 17 363 26
rect 371 17 373 26
rect 381 14 383 26
rect 388 14 390 26
rect 409 20 411 29
rect 422 18 424 29
rect 429 18 431 29
rect 450 22 452 31
rect 466 17 468 26
rect 476 17 478 26
rect 486 14 488 26
rect 493 14 495 26
rect 514 22 516 31
rect 524 25 526 31
rect 534 25 536 31
rect 554 20 556 29
rect 567 18 569 29
rect 574 18 576 29
rect 595 22 597 31
rect 611 17 613 26
rect 621 17 623 26
rect 631 14 633 26
rect 638 14 640 26
rect 659 20 661 29
rect 672 18 674 29
rect 679 18 681 29
rect 700 22 702 31
rect 716 17 718 26
rect 726 17 728 26
rect 736 14 738 26
rect 743 14 745 26
rect 764 22 766 31
rect 774 25 776 31
rect 784 25 786 31
rect 804 20 806 29
rect 817 18 819 29
rect 824 18 826 29
rect 845 22 847 31
rect 861 17 863 26
rect 871 17 873 26
rect 881 14 883 26
rect 888 14 890 26
rect 909 20 911 29
rect 922 18 924 29
rect 929 18 931 29
rect 950 22 952 31
rect 966 17 968 26
rect 976 17 978 26
rect 986 14 988 26
rect 993 14 995 26
<< pmos >>
rect 14 43 16 61
rect 27 50 29 71
rect 34 50 36 71
rect 54 44 56 62
rect 64 51 66 64
rect 74 51 76 64
rect 103 44 105 71
rect 119 44 121 62
rect 129 44 131 62
rect 139 44 141 71
rect 159 44 161 62
rect 169 51 171 64
rect 179 51 181 64
rect 208 44 210 71
rect 224 44 226 62
rect 234 44 236 62
rect 244 44 246 71
rect 264 43 266 61
rect 277 50 279 71
rect 284 50 286 71
rect 304 44 306 62
rect 314 51 316 64
rect 324 51 326 64
rect 353 44 355 71
rect 369 44 371 62
rect 379 44 381 62
rect 389 44 391 71
rect 409 44 411 62
rect 419 51 421 64
rect 429 51 431 64
rect 458 44 460 71
rect 474 44 476 62
rect 484 44 486 62
rect 494 44 496 71
rect 514 43 516 61
rect 527 50 529 71
rect 534 50 536 71
rect 554 44 556 62
rect 564 51 566 64
rect 574 51 576 64
rect 603 44 605 71
rect 619 44 621 62
rect 629 44 631 62
rect 639 44 641 71
rect 659 44 661 62
rect 669 51 671 64
rect 679 51 681 64
rect 708 44 710 71
rect 724 44 726 62
rect 734 44 736 62
rect 744 44 746 71
rect 764 43 766 61
rect 777 50 779 71
rect 784 50 786 71
rect 804 44 806 62
rect 814 51 816 64
rect 824 51 826 64
rect 853 44 855 71
rect 869 44 871 62
rect 879 44 881 62
rect 889 44 891 71
rect 909 44 911 62
rect 919 51 921 64
rect 929 51 931 64
rect 958 44 960 71
rect 974 44 976 62
rect 984 44 986 62
rect 994 44 996 71
<< polyct0 >>
rect 16 36 18 38
rect 56 36 58 38
rect 127 36 129 38
rect 137 37 139 39
rect 161 36 163 38
rect 232 36 234 38
rect 242 37 244 39
rect 266 36 268 38
rect 306 36 308 38
rect 377 36 379 38
rect 387 37 389 39
rect 411 36 413 38
rect 482 36 484 38
rect 492 37 494 39
rect 516 36 518 38
rect 556 36 558 38
rect 627 36 629 38
rect 637 37 639 39
rect 661 36 663 38
rect 732 36 734 38
rect 742 37 744 39
rect 766 36 768 38
rect 806 36 808 38
rect 877 36 879 38
rect 887 37 889 39
rect 911 36 913 38
rect 982 36 984 38
rect 992 37 994 39
<< polyct1 >>
rect 36 43 38 45
rect 26 36 28 38
rect 76 44 78 46
rect 90 44 92 46
rect 66 36 68 38
rect 181 44 183 46
rect 195 44 197 46
rect 106 31 108 33
rect 171 36 173 38
rect 286 43 288 45
rect 211 31 213 33
rect 276 36 278 38
rect 326 44 328 46
rect 340 44 342 46
rect 316 36 318 38
rect 431 44 433 46
rect 445 44 447 46
rect 356 31 358 33
rect 421 36 423 38
rect 536 43 538 45
rect 461 31 463 33
rect 526 36 528 38
rect 576 44 578 46
rect 590 44 592 46
rect 566 36 568 38
rect 681 44 683 46
rect 695 44 697 46
rect 606 31 608 33
rect 671 36 673 38
rect 786 43 788 45
rect 711 31 713 33
rect 776 36 778 38
rect 826 44 828 46
rect 840 44 842 46
rect 816 36 818 38
rect 931 44 933 46
rect 945 44 947 46
rect 856 31 858 33
rect 921 36 923 38
rect 961 31 963 33
<< ndifct0 >>
rect 29 27 31 29
rect 20 14 22 16
rect 90 27 92 29
rect 79 20 81 22
rect 104 19 106 21
rect 39 14 41 16
rect 116 22 118 24
rect 195 27 197 29
rect 184 20 186 22
rect 209 19 211 21
rect 221 22 223 24
rect 279 27 281 29
rect 270 14 272 16
rect 340 27 342 29
rect 329 20 331 22
rect 354 19 356 21
rect 289 14 291 16
rect 366 22 368 24
rect 445 27 447 29
rect 434 20 436 22
rect 459 19 461 21
rect 471 22 473 24
rect 529 27 531 29
rect 520 14 522 16
rect 590 27 592 29
rect 579 20 581 22
rect 604 19 606 21
rect 539 14 541 16
rect 616 22 618 24
rect 695 27 697 29
rect 684 20 686 22
rect 709 19 711 21
rect 721 22 723 24
rect 779 27 781 29
rect 770 14 772 16
rect 840 27 842 29
rect 829 20 831 22
rect 854 19 856 21
rect 789 14 791 16
rect 866 22 868 24
rect 945 27 947 29
rect 934 20 936 22
rect 959 19 961 21
rect 971 22 973 24
<< ndifct1 >>
rect 9 27 11 29
rect 49 22 51 24
rect 126 20 128 22
rect 60 10 62 12
rect 154 22 156 24
rect 259 27 261 29
rect 144 10 146 12
rect 231 20 233 22
rect 165 10 167 12
rect 299 22 301 24
rect 249 10 251 12
rect 376 20 378 22
rect 310 10 312 12
rect 404 22 406 24
rect 509 27 511 29
rect 394 10 396 12
rect 481 20 483 22
rect 415 10 417 12
rect 549 22 551 24
rect 499 10 501 12
rect 626 20 628 22
rect 560 10 562 12
rect 654 22 656 24
rect 759 27 761 29
rect 644 10 646 12
rect 731 20 733 22
rect 665 10 667 12
rect 799 22 801 24
rect 749 10 751 12
rect 876 20 878 22
rect 810 10 812 12
rect 904 22 906 24
rect 894 10 896 12
rect 981 20 983 22
rect 915 10 917 12
rect 999 10 1001 12
<< ntiect1 >>
rect 10 70 12 72
rect 50 70 52 72
rect 124 70 126 72
rect 155 70 157 72
rect 229 70 231 72
rect 260 70 262 72
rect 300 70 302 72
rect 374 70 376 72
rect 405 70 407 72
rect 479 70 481 72
rect 510 70 512 72
rect 550 70 552 72
rect 624 70 626 72
rect 655 70 657 72
rect 729 70 731 72
rect 760 70 762 72
rect 800 70 802 72
rect 874 70 876 72
rect 905 70 907 72
rect 979 70 981 72
<< ptiect1 >>
rect 10 10 12 12
rect 50 10 52 12
rect 91 10 93 12
rect 155 10 157 12
rect 196 10 198 12
rect 260 10 262 12
rect 300 10 302 12
rect 341 10 343 12
rect 405 10 407 12
rect 446 10 448 12
rect 510 10 512 12
rect 550 10 552 12
rect 591 10 593 12
rect 655 10 657 12
rect 696 10 698 12
rect 760 10 762 12
rect 800 10 802 12
rect 841 10 843 12
rect 905 10 907 12
rect 946 10 948 12
<< pdifct0 >>
rect 20 67 22 69
rect 39 60 41 62
rect 59 58 61 60
rect 69 60 71 62
rect 69 53 71 55
rect 79 60 81 62
rect 98 46 100 48
rect 108 67 110 69
rect 108 60 110 62
rect 124 53 126 55
rect 124 46 126 48
rect 144 61 146 63
rect 164 58 166 60
rect 174 60 176 62
rect 174 53 176 55
rect 184 60 186 62
rect 203 46 205 48
rect 213 67 215 69
rect 213 60 215 62
rect 229 53 231 55
rect 229 46 231 48
rect 270 67 272 69
rect 249 61 251 63
rect 289 60 291 62
rect 309 58 311 60
rect 319 60 321 62
rect 319 53 321 55
rect 329 60 331 62
rect 348 46 350 48
rect 358 67 360 69
rect 358 60 360 62
rect 374 53 376 55
rect 374 46 376 48
rect 394 61 396 63
rect 414 58 416 60
rect 424 60 426 62
rect 424 53 426 55
rect 434 60 436 62
rect 453 46 455 48
rect 463 67 465 69
rect 463 60 465 62
rect 479 53 481 55
rect 479 46 481 48
rect 520 67 522 69
rect 499 61 501 63
rect 539 60 541 62
rect 559 58 561 60
rect 569 60 571 62
rect 569 53 571 55
rect 579 60 581 62
rect 598 46 600 48
rect 608 67 610 69
rect 608 60 610 62
rect 624 53 626 55
rect 624 46 626 48
rect 644 61 646 63
rect 664 58 666 60
rect 674 60 676 62
rect 674 53 676 55
rect 684 60 686 62
rect 703 46 705 48
rect 713 67 715 69
rect 713 60 715 62
rect 729 53 731 55
rect 729 46 731 48
rect 770 67 772 69
rect 749 61 751 63
rect 789 60 791 62
rect 809 58 811 60
rect 819 60 821 62
rect 819 53 821 55
rect 829 60 831 62
rect 848 46 850 48
rect 858 67 860 69
rect 858 60 860 62
rect 874 53 876 55
rect 874 46 876 48
rect 894 61 896 63
rect 914 58 916 60
rect 924 60 926 62
rect 924 53 926 55
rect 934 60 936 62
rect 953 46 955 48
rect 963 67 965 69
rect 963 60 965 62
rect 979 53 981 55
rect 979 46 981 48
rect 999 61 1001 63
<< pdifct1 >>
rect 9 57 11 59
rect 9 50 11 52
rect 49 53 51 55
rect 49 46 51 48
rect 134 53 136 55
rect 154 53 156 55
rect 154 46 156 48
rect 239 53 241 55
rect 259 57 261 59
rect 259 50 261 52
rect 299 53 301 55
rect 299 46 301 48
rect 384 53 386 55
rect 404 53 406 55
rect 404 46 406 48
rect 489 53 491 55
rect 509 57 511 59
rect 509 50 511 52
rect 549 53 551 55
rect 549 46 551 48
rect 634 53 636 55
rect 654 53 656 55
rect 654 46 656 48
rect 739 53 741 55
rect 759 57 761 59
rect 759 50 761 52
rect 799 53 801 55
rect 799 46 801 48
rect 884 53 886 55
rect 904 53 906 55
rect 904 46 906 48
rect 989 53 991 55
<< alu0 >>
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 26 62 43 63
rect 26 60 39 62
rect 41 60 43 62
rect 26 59 43 60
rect 57 60 63 69
rect 11 48 12 59
rect 26 55 30 59
rect 57 58 59 60
rect 61 58 63 60
rect 57 57 63 58
rect 68 62 72 64
rect 68 60 69 62
rect 71 60 72 62
rect 15 51 30 55
rect 15 38 19 51
rect 68 55 72 60
rect 77 62 83 69
rect 107 67 108 69
rect 110 67 111 69
rect 77 60 79 62
rect 81 60 83 62
rect 77 59 83 60
rect 107 62 111 67
rect 107 60 108 62
rect 110 60 111 62
rect 107 58 111 60
rect 115 63 148 64
rect 115 61 144 63
rect 146 61 148 63
rect 115 60 148 61
rect 162 60 168 69
rect 68 54 69 55
rect 55 53 69 54
rect 71 53 72 55
rect 55 50 72 53
rect 34 42 40 43
rect 15 36 16 38
rect 18 36 19 38
rect 15 30 19 36
rect 15 29 33 30
rect 15 27 29 29
rect 31 27 33 29
rect 15 26 33 27
rect 55 38 59 50
rect 115 49 119 60
rect 162 58 164 60
rect 166 58 168 60
rect 162 57 168 58
rect 173 62 177 64
rect 173 60 174 62
rect 176 60 177 62
rect 96 48 119 49
rect 96 46 98 48
rect 100 46 119 48
rect 96 45 119 46
rect 96 39 100 45
rect 55 36 56 38
rect 58 36 59 38
rect 55 31 59 36
rect 55 27 67 31
rect 51 24 52 26
rect 63 23 67 27
rect 89 35 100 39
rect 89 29 93 35
rect 115 39 119 45
rect 123 55 127 57
rect 123 53 124 55
rect 126 53 127 55
rect 123 48 127 53
rect 123 46 124 48
rect 126 47 127 48
rect 126 46 139 47
rect 123 43 139 46
rect 135 41 139 43
rect 135 39 140 41
rect 115 38 131 39
rect 115 36 127 38
rect 129 36 131 38
rect 115 35 131 36
rect 135 37 137 39
rect 139 37 140 39
rect 135 35 140 37
rect 89 27 90 29
rect 92 27 93 29
rect 89 25 93 27
rect 135 31 139 35
rect 115 27 139 31
rect 115 24 119 27
rect 63 22 83 23
rect 115 22 116 24
rect 118 22 119 24
rect 63 20 79 22
rect 81 20 83 22
rect 63 19 83 20
rect 102 21 108 22
rect 102 19 104 21
rect 106 19 108 21
rect 115 20 119 22
rect 173 55 177 60
rect 182 62 188 69
rect 212 67 213 69
rect 215 67 216 69
rect 182 60 184 62
rect 186 60 188 62
rect 182 59 188 60
rect 212 62 216 67
rect 268 67 270 69
rect 272 67 274 69
rect 268 66 274 67
rect 212 60 213 62
rect 215 60 216 62
rect 212 58 216 60
rect 220 63 253 64
rect 220 61 249 63
rect 251 61 253 63
rect 220 60 253 61
rect 173 54 174 55
rect 160 53 174 54
rect 176 53 177 55
rect 160 50 177 53
rect 160 38 164 50
rect 220 49 224 60
rect 276 62 293 63
rect 276 60 289 62
rect 291 60 293 62
rect 276 59 293 60
rect 307 60 313 69
rect 201 48 224 49
rect 201 46 203 48
rect 205 46 224 48
rect 201 45 224 46
rect 201 39 205 45
rect 160 36 161 38
rect 163 36 164 38
rect 160 31 164 36
rect 160 27 172 31
rect 156 24 157 26
rect 18 16 24 17
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 37 16 43 17
rect 37 14 39 16
rect 41 14 43 16
rect 37 13 43 14
rect 102 13 108 19
rect 168 23 172 27
rect 194 35 205 39
rect 194 29 198 35
rect 220 39 224 45
rect 228 55 232 57
rect 228 53 229 55
rect 231 53 232 55
rect 228 48 232 53
rect 228 46 229 48
rect 231 47 232 48
rect 231 46 244 47
rect 228 43 244 46
rect 240 41 244 43
rect 240 39 245 41
rect 220 38 236 39
rect 220 36 232 38
rect 234 36 236 38
rect 220 35 236 36
rect 240 37 242 39
rect 244 37 245 39
rect 240 35 245 37
rect 194 27 195 29
rect 197 27 198 29
rect 194 25 198 27
rect 240 31 244 35
rect 220 27 244 31
rect 220 24 224 27
rect 168 22 188 23
rect 220 22 221 24
rect 223 22 224 24
rect 261 48 262 59
rect 276 55 280 59
rect 307 58 309 60
rect 311 58 313 60
rect 307 57 313 58
rect 318 62 322 64
rect 318 60 319 62
rect 321 60 322 62
rect 265 51 280 55
rect 265 38 269 51
rect 318 55 322 60
rect 327 62 333 69
rect 357 67 358 69
rect 360 67 361 69
rect 327 60 329 62
rect 331 60 333 62
rect 327 59 333 60
rect 357 62 361 67
rect 357 60 358 62
rect 360 60 361 62
rect 357 58 361 60
rect 365 63 398 64
rect 365 61 394 63
rect 396 61 398 63
rect 365 60 398 61
rect 412 60 418 69
rect 318 54 319 55
rect 305 53 319 54
rect 321 53 322 55
rect 305 50 322 53
rect 284 42 290 43
rect 265 36 266 38
rect 268 36 269 38
rect 265 30 269 36
rect 265 29 283 30
rect 265 27 279 29
rect 281 27 283 29
rect 265 26 283 27
rect 168 20 184 22
rect 186 20 188 22
rect 168 19 188 20
rect 207 21 213 22
rect 207 19 209 21
rect 211 19 213 21
rect 220 20 224 22
rect 305 38 309 50
rect 365 49 369 60
rect 412 58 414 60
rect 416 58 418 60
rect 412 57 418 58
rect 423 62 427 64
rect 423 60 424 62
rect 426 60 427 62
rect 346 48 369 49
rect 346 46 348 48
rect 350 46 369 48
rect 346 45 369 46
rect 346 39 350 45
rect 305 36 306 38
rect 308 36 309 38
rect 305 31 309 36
rect 305 27 317 31
rect 301 24 302 26
rect 207 13 213 19
rect 313 23 317 27
rect 339 35 350 39
rect 339 29 343 35
rect 365 39 369 45
rect 373 55 377 57
rect 373 53 374 55
rect 376 53 377 55
rect 373 48 377 53
rect 373 46 374 48
rect 376 47 377 48
rect 376 46 389 47
rect 373 43 389 46
rect 385 41 389 43
rect 385 39 390 41
rect 365 38 381 39
rect 365 36 377 38
rect 379 36 381 38
rect 365 35 381 36
rect 385 37 387 39
rect 389 37 390 39
rect 385 35 390 37
rect 339 27 340 29
rect 342 27 343 29
rect 339 25 343 27
rect 385 31 389 35
rect 365 27 389 31
rect 365 24 369 27
rect 313 22 333 23
rect 365 22 366 24
rect 368 22 369 24
rect 313 20 329 22
rect 331 20 333 22
rect 313 19 333 20
rect 352 21 358 22
rect 352 19 354 21
rect 356 19 358 21
rect 365 20 369 22
rect 423 55 427 60
rect 432 62 438 69
rect 462 67 463 69
rect 465 67 466 69
rect 432 60 434 62
rect 436 60 438 62
rect 432 59 438 60
rect 462 62 466 67
rect 518 67 520 69
rect 522 67 524 69
rect 518 66 524 67
rect 462 60 463 62
rect 465 60 466 62
rect 462 58 466 60
rect 470 63 503 64
rect 470 61 499 63
rect 501 61 503 63
rect 470 60 503 61
rect 423 54 424 55
rect 410 53 424 54
rect 426 53 427 55
rect 410 50 427 53
rect 410 38 414 50
rect 470 49 474 60
rect 526 62 543 63
rect 526 60 539 62
rect 541 60 543 62
rect 526 59 543 60
rect 557 60 563 69
rect 451 48 474 49
rect 451 46 453 48
rect 455 46 474 48
rect 451 45 474 46
rect 451 39 455 45
rect 410 36 411 38
rect 413 36 414 38
rect 410 31 414 36
rect 410 27 422 31
rect 406 24 407 26
rect 268 16 274 17
rect 268 14 270 16
rect 272 14 274 16
rect 268 13 274 14
rect 287 16 293 17
rect 287 14 289 16
rect 291 14 293 16
rect 287 13 293 14
rect 352 13 358 19
rect 418 23 422 27
rect 444 35 455 39
rect 444 29 448 35
rect 470 39 474 45
rect 478 55 482 57
rect 478 53 479 55
rect 481 53 482 55
rect 478 48 482 53
rect 478 46 479 48
rect 481 47 482 48
rect 481 46 494 47
rect 478 43 494 46
rect 490 41 494 43
rect 490 39 495 41
rect 470 38 486 39
rect 470 36 482 38
rect 484 36 486 38
rect 470 35 486 36
rect 490 37 492 39
rect 494 37 495 39
rect 490 35 495 37
rect 444 27 445 29
rect 447 27 448 29
rect 444 25 448 27
rect 490 31 494 35
rect 470 27 494 31
rect 470 24 474 27
rect 418 22 438 23
rect 470 22 471 24
rect 473 22 474 24
rect 511 48 512 59
rect 526 55 530 59
rect 557 58 559 60
rect 561 58 563 60
rect 557 57 563 58
rect 568 62 572 64
rect 568 60 569 62
rect 571 60 572 62
rect 515 51 530 55
rect 515 38 519 51
rect 568 55 572 60
rect 577 62 583 69
rect 607 67 608 69
rect 610 67 611 69
rect 577 60 579 62
rect 581 60 583 62
rect 577 59 583 60
rect 607 62 611 67
rect 607 60 608 62
rect 610 60 611 62
rect 607 58 611 60
rect 615 63 648 64
rect 615 61 644 63
rect 646 61 648 63
rect 615 60 648 61
rect 662 60 668 69
rect 568 54 569 55
rect 555 53 569 54
rect 571 53 572 55
rect 555 50 572 53
rect 534 42 540 43
rect 515 36 516 38
rect 518 36 519 38
rect 515 30 519 36
rect 515 29 533 30
rect 515 27 529 29
rect 531 27 533 29
rect 515 26 533 27
rect 418 20 434 22
rect 436 20 438 22
rect 418 19 438 20
rect 457 21 463 22
rect 457 19 459 21
rect 461 19 463 21
rect 470 20 474 22
rect 555 38 559 50
rect 615 49 619 60
rect 662 58 664 60
rect 666 58 668 60
rect 662 57 668 58
rect 673 62 677 64
rect 673 60 674 62
rect 676 60 677 62
rect 596 48 619 49
rect 596 46 598 48
rect 600 46 619 48
rect 596 45 619 46
rect 596 39 600 45
rect 555 36 556 38
rect 558 36 559 38
rect 555 31 559 36
rect 555 27 567 31
rect 551 24 552 26
rect 457 13 463 19
rect 563 23 567 27
rect 589 35 600 39
rect 589 29 593 35
rect 615 39 619 45
rect 623 55 627 57
rect 623 53 624 55
rect 626 53 627 55
rect 623 48 627 53
rect 623 46 624 48
rect 626 47 627 48
rect 626 46 639 47
rect 623 43 639 46
rect 635 41 639 43
rect 635 39 640 41
rect 615 38 631 39
rect 615 36 627 38
rect 629 36 631 38
rect 615 35 631 36
rect 635 37 637 39
rect 639 37 640 39
rect 635 35 640 37
rect 589 27 590 29
rect 592 27 593 29
rect 589 25 593 27
rect 635 31 639 35
rect 615 27 639 31
rect 615 24 619 27
rect 563 22 583 23
rect 615 22 616 24
rect 618 22 619 24
rect 563 20 579 22
rect 581 20 583 22
rect 563 19 583 20
rect 602 21 608 22
rect 602 19 604 21
rect 606 19 608 21
rect 615 20 619 22
rect 673 55 677 60
rect 682 62 688 69
rect 712 67 713 69
rect 715 67 716 69
rect 682 60 684 62
rect 686 60 688 62
rect 682 59 688 60
rect 712 62 716 67
rect 768 67 770 69
rect 772 67 774 69
rect 768 66 774 67
rect 712 60 713 62
rect 715 60 716 62
rect 712 58 716 60
rect 720 63 753 64
rect 720 61 749 63
rect 751 61 753 63
rect 720 60 753 61
rect 673 54 674 55
rect 660 53 674 54
rect 676 53 677 55
rect 660 50 677 53
rect 660 38 664 50
rect 720 49 724 60
rect 776 62 793 63
rect 776 60 789 62
rect 791 60 793 62
rect 776 59 793 60
rect 807 60 813 69
rect 701 48 724 49
rect 701 46 703 48
rect 705 46 724 48
rect 701 45 724 46
rect 701 39 705 45
rect 660 36 661 38
rect 663 36 664 38
rect 660 31 664 36
rect 660 27 672 31
rect 656 24 657 26
rect 518 16 524 17
rect 518 14 520 16
rect 522 14 524 16
rect 518 13 524 14
rect 537 16 543 17
rect 537 14 539 16
rect 541 14 543 16
rect 537 13 543 14
rect 602 13 608 19
rect 668 23 672 27
rect 694 35 705 39
rect 694 29 698 35
rect 720 39 724 45
rect 728 55 732 57
rect 728 53 729 55
rect 731 53 732 55
rect 728 48 732 53
rect 728 46 729 48
rect 731 47 732 48
rect 731 46 744 47
rect 728 43 744 46
rect 740 41 744 43
rect 740 39 745 41
rect 720 38 736 39
rect 720 36 732 38
rect 734 36 736 38
rect 720 35 736 36
rect 740 37 742 39
rect 744 37 745 39
rect 740 35 745 37
rect 694 27 695 29
rect 697 27 698 29
rect 694 25 698 27
rect 740 31 744 35
rect 720 27 744 31
rect 720 24 724 27
rect 668 22 688 23
rect 720 22 721 24
rect 723 22 724 24
rect 761 48 762 59
rect 776 55 780 59
rect 807 58 809 60
rect 811 58 813 60
rect 807 57 813 58
rect 818 62 822 64
rect 818 60 819 62
rect 821 60 822 62
rect 765 51 780 55
rect 765 38 769 51
rect 818 55 822 60
rect 827 62 833 69
rect 857 67 858 69
rect 860 67 861 69
rect 827 60 829 62
rect 831 60 833 62
rect 827 59 833 60
rect 857 62 861 67
rect 857 60 858 62
rect 860 60 861 62
rect 857 58 861 60
rect 865 63 898 64
rect 865 61 894 63
rect 896 61 898 63
rect 865 60 898 61
rect 912 60 918 69
rect 818 54 819 55
rect 805 53 819 54
rect 821 53 822 55
rect 805 50 822 53
rect 784 42 790 43
rect 765 36 766 38
rect 768 36 769 38
rect 765 30 769 36
rect 765 29 783 30
rect 765 27 779 29
rect 781 27 783 29
rect 765 26 783 27
rect 668 20 684 22
rect 686 20 688 22
rect 668 19 688 20
rect 707 21 713 22
rect 707 19 709 21
rect 711 19 713 21
rect 720 20 724 22
rect 805 38 809 50
rect 865 49 869 60
rect 912 58 914 60
rect 916 58 918 60
rect 912 57 918 58
rect 923 62 927 64
rect 923 60 924 62
rect 926 60 927 62
rect 846 48 869 49
rect 846 46 848 48
rect 850 46 869 48
rect 846 45 869 46
rect 846 39 850 45
rect 805 36 806 38
rect 808 36 809 38
rect 805 31 809 36
rect 805 27 817 31
rect 801 24 802 26
rect 707 13 713 19
rect 813 23 817 27
rect 839 35 850 39
rect 839 29 843 35
rect 865 39 869 45
rect 873 55 877 57
rect 873 53 874 55
rect 876 53 877 55
rect 873 48 877 53
rect 873 46 874 48
rect 876 47 877 48
rect 876 46 889 47
rect 873 43 889 46
rect 885 41 889 43
rect 885 39 890 41
rect 865 38 881 39
rect 865 36 877 38
rect 879 36 881 38
rect 865 35 881 36
rect 885 37 887 39
rect 889 37 890 39
rect 885 35 890 37
rect 839 27 840 29
rect 842 27 843 29
rect 839 25 843 27
rect 885 31 889 35
rect 865 27 889 31
rect 865 24 869 27
rect 813 22 833 23
rect 865 22 866 24
rect 868 22 869 24
rect 813 20 829 22
rect 831 20 833 22
rect 813 19 833 20
rect 852 21 858 22
rect 852 19 854 21
rect 856 19 858 21
rect 865 20 869 22
rect 923 55 927 60
rect 932 62 938 69
rect 962 67 963 69
rect 965 67 966 69
rect 932 60 934 62
rect 936 60 938 62
rect 932 59 938 60
rect 962 62 966 67
rect 962 60 963 62
rect 965 60 966 62
rect 962 58 966 60
rect 970 63 1003 64
rect 970 61 999 63
rect 1001 61 1003 63
rect 970 60 1003 61
rect 923 54 924 55
rect 910 53 924 54
rect 926 53 927 55
rect 910 50 927 53
rect 910 38 914 50
rect 970 49 974 60
rect 951 48 974 49
rect 951 46 953 48
rect 955 46 974 48
rect 951 45 974 46
rect 951 39 955 45
rect 910 36 911 38
rect 913 36 914 38
rect 910 31 914 36
rect 910 27 922 31
rect 906 24 907 26
rect 768 16 774 17
rect 768 14 770 16
rect 772 14 774 16
rect 768 13 774 14
rect 787 16 793 17
rect 787 14 789 16
rect 791 14 793 16
rect 787 13 793 14
rect 852 13 858 19
rect 918 23 922 27
rect 944 35 955 39
rect 944 29 948 35
rect 970 39 974 45
rect 978 55 982 57
rect 978 53 979 55
rect 981 53 982 55
rect 978 48 982 53
rect 978 46 979 48
rect 981 47 982 48
rect 981 46 994 47
rect 978 43 994 46
rect 990 41 994 43
rect 990 39 995 41
rect 970 38 986 39
rect 970 36 982 38
rect 984 36 986 38
rect 970 35 986 36
rect 990 37 992 39
rect 994 37 995 39
rect 990 35 995 37
rect 944 27 945 29
rect 947 27 948 29
rect 944 25 948 27
rect 990 31 994 35
rect 970 27 994 31
rect 970 24 974 27
rect 918 22 938 23
rect 970 22 971 24
rect 973 22 974 24
rect 918 20 934 22
rect 936 20 938 22
rect 918 19 938 20
rect 957 21 963 22
rect 957 19 959 21
rect 961 19 963 21
rect 970 20 974 22
rect 957 13 963 19
<< via1 >>
rect 40 53 42 55
rect 72 27 74 29
rect 99 27 101 29
rect 145 27 147 29
rect 154 53 156 55
rect 187 45 189 47
rect 177 27 179 29
rect 204 27 206 29
rect 290 53 292 55
rect 258 45 260 47
rect 322 27 324 29
rect 349 27 351 29
rect 395 27 397 29
rect 404 53 406 55
rect 439 45 441 47
rect 427 27 429 29
rect 454 27 456 29
rect 540 53 542 55
rect 508 45 510 47
rect 572 27 574 29
rect 599 27 601 29
rect 645 27 647 29
rect 654 53 656 55
rect 689 45 691 47
rect 677 27 679 29
rect 704 27 706 29
rect 790 53 792 55
rect 758 45 760 47
rect 822 27 824 29
rect 849 27 851 29
rect 895 27 897 29
rect 904 53 906 55
rect 939 44 941 46
rect 927 27 929 29
rect 954 27 956 29
rect 939 9 941 11
<< via2 >>
rect 939 35 941 37
rect 939 19 941 21
<< labels >>
rlabel alu1 89 73 89 73 1 Vdd
rlabel alu1 65 73 65 73 6 vdd
rlabel alu1 87 8 87 8 1 Vss
rlabel alu1 194 73 194 73 1 Vdd
rlabel alu1 170 73 170 73 6 vdd
rlabel alu1 192 8 192 8 1 Vss
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 339 73 339 73 1 Vdd
rlabel alu1 315 73 315 73 6 vdd
rlabel alu1 337 8 337 8 1 Vss
rlabel alu1 444 73 444 73 1 Vdd
rlabel alu1 420 73 420 73 6 vdd
rlabel alu1 442 8 442 8 1 Vss
rlabel alu1 275 73 275 73 6 vdd
rlabel alu1 525 73 525 73 6 vdd
rlabel alu1 692 8 692 8 1 Vss
rlabel alu1 670 73 670 73 6 vdd
rlabel alu1 694 73 694 73 1 Vdd
rlabel alu1 587 8 587 8 1 Vss
rlabel alu1 565 73 565 73 6 vdd
rlabel alu1 589 73 589 73 1 Vdd
rlabel alu1 839 73 839 73 1 Vdd
rlabel alu1 815 73 815 73 6 vdd
rlabel alu1 837 8 837 8 1 Vss
rlabel alu1 944 73 944 73 1 Vdd
rlabel alu1 920 73 920 73 6 vdd
rlabel alu1 942 8 942 8 1 Vss
rlabel alu1 775 73 775 73 6 vdd
rlabel alu1 936 53 936 53 1 Vss
rlabel alu1 9 44 9 44 1 c2
rlabel alu1 98 61 98 61 1 p33
rlabel alu1 348 61 348 61 1 p32
rlabel alu1 598 61 598 61 1 p31
rlabel alu1 607 36 607 36 1 s13
rlabel alu1 848 61 848 61 1 p30
rlabel alu1 857 36 857 36 1 s12
rlabel alu1 1001 40 1001 40 1 r4
rlabel alu1 751 40 751 40 1 r5
rlabel alu1 501 40 501 40 1 r6
rlabel alu1 251 40 251 40 1 r7
rlabel alu1 357 36 357 36 1 sha
rlabel alu1 107 36 107 36 1 cha
<< end >>
