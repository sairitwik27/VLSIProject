magic
tech scmos
timestamp 1609005231
<< ab >>
rect 23 223 71 231
rect 32 158 71 223
rect 73 158 109 231
rect 32 95 69 158
rect 23 91 69 95
rect 71 91 109 158
rect 23 87 109 91
rect 111 223 116 231
rect 111 167 113 223
rect 111 158 116 167
rect 118 158 181 231
rect 183 199 221 231
rect 353 222 399 229
rect 183 158 230 199
rect 362 159 399 222
rect 401 159 439 229
rect 111 87 151 158
rect 153 87 216 158
rect 221 119 230 158
rect 235 95 275 159
rect 217 87 275 95
rect 277 87 340 159
rect 362 94 401 159
rect 341 87 401 94
rect 353 86 401 87
rect 403 87 439 159
rect 441 159 481 229
rect 483 159 546 229
rect 548 222 604 229
rect 551 166 560 198
rect 567 166 604 222
rect 551 159 604 166
rect 606 159 644 229
rect 441 150 446 159
rect 441 94 443 150
rect 441 87 446 94
rect 403 86 446 87
rect 448 86 511 159
rect 513 150 606 159
rect 513 118 560 150
rect 513 94 551 118
rect 567 94 606 150
rect 513 86 606 94
rect 608 86 644 159
rect 646 159 686 229
rect 688 159 751 229
rect 1813 223 1861 231
rect 756 159 765 198
rect 646 150 651 159
rect 646 94 648 150
rect 646 86 651 94
rect 653 86 716 159
rect 718 118 765 159
rect 718 86 756 118
rect 773 87 853 159
rect 855 87 958 159
rect 960 87 1103 159
rect 1105 87 1208 159
rect 1210 87 1353 159
rect 1355 87 1458 159
rect 1460 87 1603 159
rect 1605 87 1708 159
rect 1710 87 1773 159
rect 1822 158 1861 223
rect 1863 158 1899 231
rect 1775 151 1859 158
rect 1822 95 1859 151
rect 1775 88 1859 95
rect 1813 87 1859 88
rect 1861 87 1899 158
rect 1901 223 1906 231
rect 1901 167 1903 223
rect 1901 158 1906 167
rect 1908 158 1971 231
rect 1973 199 2011 231
rect 1973 158 2020 199
rect 1901 87 1941 158
rect 1943 87 2006 158
rect 2011 119 2020 158
rect 1031 86 1077 87
rect 1079 86 1117 87
rect 1119 86 1159 87
rect 1161 86 1224 87
rect 1226 86 1282 87
rect 1284 86 1322 87
rect 1324 86 1364 87
rect 1366 86 1429 87
rect 436 77 441 86
rect 5 5 85 77
rect 87 69 190 77
rect 87 60 100 69
rect 102 60 190 69
rect 87 5 190 60
rect 192 5 335 77
rect 337 5 440 77
rect 442 5 585 77
rect 587 5 690 77
rect 692 5 835 77
rect 837 50 940 77
rect 942 50 1005 77
rect 837 48 1005 50
rect 837 5 940 48
rect 942 5 1005 48
rect 1015 13 1095 77
rect 1007 5 1095 13
rect 1097 5 1200 77
rect 1202 39 1345 77
rect 1347 39 1450 77
rect 1202 38 1450 39
rect 1202 5 1345 38
rect 1347 5 1450 38
rect 1452 39 1595 77
rect 1597 39 1700 77
rect 1452 37 1700 39
rect 1452 5 1595 37
rect 1597 5 1700 37
rect 1702 5 1845 77
rect 1847 50 1950 77
rect 1952 50 2015 77
rect 1847 48 2015 50
rect 1847 5 1950 48
rect 1952 5 2015 48
<< nwell >>
rect 14 198 230 199
rect 1804 198 2020 199
rect 14 119 2020 198
rect 344 118 767 119
rect 1778 118 1804 119
rect 0 0 2020 45
<< pwell >>
rect 345 236 766 237
rect 14 199 2020 236
rect 230 198 1804 199
rect 14 118 344 119
rect 767 118 1778 119
rect 1804 118 2020 119
rect 14 82 2020 118
rect 0 45 2020 82
<< poly >>
rect 40 218 42 223
rect 47 218 49 223
rect 60 216 62 220
rect 80 218 82 223
rect 87 218 89 223
rect 145 227 170 229
rect 128 222 130 227
rect 135 222 137 227
rect 100 216 102 220
rect 145 219 147 227
rect 155 219 157 223
rect 168 219 170 227
rect 168 217 173 219
rect 192 218 194 223
rect 199 218 201 223
rect 171 214 173 217
rect 40 194 42 207
rect 47 202 49 207
rect 60 202 62 207
rect 46 200 52 202
rect 46 198 48 200
rect 50 198 52 200
rect 46 196 52 198
rect 56 200 62 202
rect 56 198 58 200
rect 60 198 62 200
rect 56 196 62 198
rect 36 192 42 194
rect 36 190 38 192
rect 40 190 42 192
rect 36 188 42 190
rect 40 185 42 188
rect 50 185 52 196
rect 60 192 62 196
rect 80 194 82 207
rect 87 202 89 207
rect 100 202 102 207
rect 86 200 92 202
rect 86 198 88 200
rect 90 198 92 200
rect 86 196 92 198
rect 96 200 102 202
rect 128 201 130 210
rect 135 207 137 210
rect 135 205 139 207
rect 145 206 147 210
rect 155 207 157 210
rect 137 202 139 205
rect 155 205 164 207
rect 212 216 214 220
rect 370 215 372 219
rect 383 217 385 222
rect 390 217 392 222
rect 410 217 412 222
rect 417 217 419 222
rect 155 203 160 205
rect 162 203 164 205
rect 96 198 98 200
rect 100 198 102 200
rect 96 196 102 198
rect 76 192 82 194
rect 76 190 78 192
rect 80 190 82 192
rect 76 188 82 190
rect 80 185 82 188
rect 90 185 92 196
rect 100 192 102 196
rect 127 199 133 201
rect 127 197 129 199
rect 131 197 133 199
rect 127 195 133 197
rect 137 200 143 202
rect 137 198 139 200
rect 141 198 143 200
rect 137 196 143 198
rect 155 201 164 203
rect 155 197 157 201
rect 171 197 173 205
rect 127 192 129 195
rect 137 192 139 196
rect 147 195 157 197
rect 163 195 176 197
rect 147 192 149 195
rect 163 192 165 195
rect 174 194 176 195
rect 192 194 194 207
rect 199 202 201 207
rect 212 202 214 207
rect 430 215 432 219
rect 450 215 452 219
rect 463 217 465 222
rect 470 217 472 222
rect 494 226 519 228
rect 494 218 496 226
rect 507 218 509 222
rect 517 218 519 226
rect 527 221 529 226
rect 534 221 536 226
rect 491 216 496 218
rect 491 213 493 216
rect 198 200 204 202
rect 198 198 200 200
rect 202 198 204 200
rect 198 196 204 198
rect 208 200 214 202
rect 208 198 210 200
rect 212 198 214 200
rect 208 196 214 198
rect 174 192 180 194
rect 40 167 42 172
rect 50 167 52 172
rect 60 170 62 174
rect 80 167 82 172
rect 90 167 92 172
rect 100 170 102 174
rect 137 170 139 174
rect 147 170 149 174
rect 127 161 129 165
rect 174 190 176 192
rect 178 190 180 192
rect 174 188 180 190
rect 188 192 194 194
rect 188 190 190 192
rect 192 190 194 192
rect 188 188 194 190
rect 192 185 194 188
rect 202 185 204 196
rect 212 192 214 196
rect 370 201 372 206
rect 383 201 385 206
rect 370 199 376 201
rect 370 197 372 199
rect 374 197 376 199
rect 370 195 376 197
rect 380 199 386 201
rect 380 197 382 199
rect 384 197 386 199
rect 380 195 386 197
rect 370 191 372 195
rect 192 167 194 172
rect 202 167 204 172
rect 212 170 214 174
rect 380 184 382 195
rect 390 193 392 206
rect 410 193 412 206
rect 417 201 419 206
rect 430 201 432 206
rect 416 199 422 201
rect 416 197 418 199
rect 420 197 422 199
rect 416 195 422 197
rect 426 199 432 201
rect 426 197 428 199
rect 430 197 432 199
rect 426 195 432 197
rect 390 191 396 193
rect 390 189 392 191
rect 394 189 396 191
rect 390 187 396 189
rect 406 191 412 193
rect 406 189 408 191
rect 410 189 412 191
rect 406 187 412 189
rect 390 184 392 187
rect 410 184 412 187
rect 420 184 422 195
rect 430 191 432 195
rect 450 201 452 206
rect 463 201 465 206
rect 450 199 456 201
rect 450 197 452 199
rect 454 197 456 199
rect 450 195 456 197
rect 460 199 466 201
rect 460 197 462 199
rect 464 197 466 199
rect 460 195 466 197
rect 450 191 452 195
rect 370 169 372 173
rect 460 184 462 195
rect 470 193 472 206
rect 575 215 577 219
rect 588 217 590 222
rect 595 217 597 222
rect 615 217 617 222
rect 622 217 624 222
rect 507 206 509 209
rect 500 204 509 206
rect 517 205 519 209
rect 527 206 529 209
rect 491 196 493 204
rect 500 202 502 204
rect 504 202 509 204
rect 500 200 509 202
rect 525 204 529 206
rect 525 201 527 204
rect 507 196 509 200
rect 521 199 527 201
rect 534 200 536 209
rect 635 215 637 219
rect 655 215 657 219
rect 668 217 670 222
rect 675 217 677 222
rect 699 226 724 228
rect 699 218 701 226
rect 712 218 714 222
rect 722 218 724 226
rect 732 221 734 226
rect 739 221 741 226
rect 696 216 701 218
rect 696 213 698 216
rect 575 201 577 206
rect 588 201 590 206
rect 521 197 523 199
rect 525 197 527 199
rect 488 194 501 196
rect 507 194 517 196
rect 521 195 527 197
rect 488 193 490 194
rect 470 191 476 193
rect 470 189 472 191
rect 474 189 476 191
rect 470 187 476 189
rect 484 191 490 193
rect 499 191 501 194
rect 515 191 517 194
rect 525 191 527 195
rect 531 198 537 200
rect 531 196 533 198
rect 535 196 537 198
rect 531 194 537 196
rect 535 191 537 194
rect 575 199 581 201
rect 575 197 577 199
rect 579 197 581 199
rect 575 195 581 197
rect 585 199 591 201
rect 585 197 587 199
rect 589 197 591 199
rect 585 195 591 197
rect 575 191 577 195
rect 484 189 486 191
rect 488 189 490 191
rect 484 187 490 189
rect 470 184 472 187
rect 163 161 165 165
rect 380 166 382 171
rect 390 166 392 171
rect 410 166 412 171
rect 420 166 422 171
rect 430 169 432 173
rect 450 169 452 173
rect 460 166 462 171
rect 470 166 472 171
rect 515 169 517 173
rect 525 169 527 173
rect 499 160 501 164
rect 585 184 587 195
rect 595 193 597 206
rect 615 193 617 206
rect 622 201 624 206
rect 635 201 637 206
rect 621 199 627 201
rect 621 197 623 199
rect 625 197 627 199
rect 621 195 627 197
rect 631 199 637 201
rect 631 197 633 199
rect 635 197 637 199
rect 631 195 637 197
rect 595 191 601 193
rect 595 189 597 191
rect 599 189 601 191
rect 595 187 601 189
rect 611 191 617 193
rect 611 189 613 191
rect 615 189 617 191
rect 611 187 617 189
rect 595 184 597 187
rect 615 184 617 187
rect 625 184 627 195
rect 635 191 637 195
rect 655 201 657 206
rect 668 201 670 206
rect 655 199 661 201
rect 655 197 657 199
rect 659 197 661 199
rect 655 195 661 197
rect 665 199 671 201
rect 665 197 667 199
rect 669 197 671 199
rect 665 195 671 197
rect 655 191 657 195
rect 575 169 577 173
rect 665 184 667 195
rect 675 193 677 206
rect 1830 218 1832 223
rect 1837 218 1839 223
rect 712 206 714 209
rect 705 204 714 206
rect 722 205 724 209
rect 732 206 734 209
rect 696 196 698 204
rect 705 202 707 204
rect 709 202 714 204
rect 705 200 714 202
rect 730 204 734 206
rect 730 201 732 204
rect 712 196 714 200
rect 726 199 732 201
rect 739 200 741 209
rect 1850 216 1852 220
rect 1870 218 1872 223
rect 1877 218 1879 223
rect 1935 227 1960 229
rect 1918 222 1920 227
rect 1925 222 1927 227
rect 1890 216 1892 220
rect 1935 219 1937 227
rect 1945 219 1947 223
rect 1958 219 1960 227
rect 1958 217 1963 219
rect 1982 218 1984 223
rect 1989 218 1991 223
rect 1961 214 1963 217
rect 726 197 728 199
rect 730 197 732 199
rect 693 194 706 196
rect 712 194 722 196
rect 726 195 732 197
rect 693 193 695 194
rect 675 191 681 193
rect 675 189 677 191
rect 679 189 681 191
rect 675 187 681 189
rect 689 191 695 193
rect 704 191 706 194
rect 720 191 722 194
rect 730 191 732 195
rect 736 198 742 200
rect 736 196 738 198
rect 740 196 742 198
rect 736 194 742 196
rect 1830 194 1832 207
rect 1837 202 1839 207
rect 1850 202 1852 207
rect 1836 200 1842 202
rect 1836 198 1838 200
rect 1840 198 1842 200
rect 1836 196 1842 198
rect 1846 200 1852 202
rect 1846 198 1848 200
rect 1850 198 1852 200
rect 1846 196 1852 198
rect 740 191 742 194
rect 1826 192 1832 194
rect 689 189 691 191
rect 693 189 695 191
rect 689 187 695 189
rect 675 184 677 187
rect 585 166 587 171
rect 595 166 597 171
rect 615 166 617 171
rect 625 166 627 171
rect 635 169 637 173
rect 655 169 657 173
rect 535 160 537 164
rect 665 166 667 171
rect 675 166 677 171
rect 720 169 722 173
rect 730 169 732 173
rect 704 160 706 164
rect 1826 190 1828 192
rect 1830 190 1832 192
rect 1826 188 1832 190
rect 1830 185 1832 188
rect 1840 185 1842 196
rect 1850 192 1852 196
rect 1870 194 1872 207
rect 1877 202 1879 207
rect 1890 202 1892 207
rect 1876 200 1882 202
rect 1876 198 1878 200
rect 1880 198 1882 200
rect 1876 196 1882 198
rect 1886 200 1892 202
rect 1918 201 1920 210
rect 1925 207 1927 210
rect 1925 205 1929 207
rect 1935 206 1937 210
rect 1945 207 1947 210
rect 1927 202 1929 205
rect 1945 205 1954 207
rect 2002 216 2004 220
rect 1945 203 1950 205
rect 1952 203 1954 205
rect 1886 198 1888 200
rect 1890 198 1892 200
rect 1886 196 1892 198
rect 1866 192 1872 194
rect 1866 190 1868 192
rect 1870 190 1872 192
rect 1866 188 1872 190
rect 1870 185 1872 188
rect 1880 185 1882 196
rect 1890 192 1892 196
rect 1917 199 1923 201
rect 1917 197 1919 199
rect 1921 197 1923 199
rect 1917 195 1923 197
rect 1927 200 1933 202
rect 1927 198 1929 200
rect 1931 198 1933 200
rect 1927 196 1933 198
rect 1945 201 1954 203
rect 1945 197 1947 201
rect 1961 197 1963 205
rect 1917 192 1919 195
rect 1927 192 1929 196
rect 1937 195 1947 197
rect 1953 195 1966 197
rect 1937 192 1939 195
rect 1953 192 1955 195
rect 1964 194 1966 195
rect 1982 194 1984 207
rect 1989 202 1991 207
rect 2002 202 2004 207
rect 1988 200 1994 202
rect 1988 198 1990 200
rect 1992 198 1994 200
rect 1988 196 1994 198
rect 1998 200 2004 202
rect 1998 198 2000 200
rect 2002 198 2004 200
rect 1998 196 2004 198
rect 1964 192 1970 194
rect 1830 167 1832 172
rect 1840 167 1842 172
rect 1850 170 1852 174
rect 1870 167 1872 172
rect 1880 167 1882 172
rect 1890 170 1892 174
rect 740 160 742 164
rect 1927 170 1929 174
rect 1937 170 1939 174
rect 1917 161 1919 165
rect 1964 190 1966 192
rect 1968 190 1970 192
rect 1964 188 1970 190
rect 1978 192 1984 194
rect 1978 190 1980 192
rect 1982 190 1984 192
rect 1978 188 1984 190
rect 1982 185 1984 188
rect 1992 185 1994 196
rect 2002 192 2004 196
rect 1982 167 1984 172
rect 1992 167 1994 172
rect 2002 170 2004 174
rect 1953 161 1955 165
rect 40 144 42 148
rect 50 146 52 151
rect 60 146 62 151
rect 80 146 82 151
rect 90 146 92 151
rect 169 153 171 157
rect 100 144 102 148
rect 120 144 122 148
rect 130 146 132 151
rect 140 146 142 151
rect 40 122 42 126
rect 50 122 52 133
rect 60 130 62 133
rect 80 130 82 133
rect 60 128 66 130
rect 60 126 62 128
rect 64 126 66 128
rect 60 124 66 126
rect 76 128 82 130
rect 76 126 78 128
rect 80 126 82 128
rect 76 124 82 126
rect 40 120 46 122
rect 40 118 42 120
rect 44 118 46 120
rect 40 116 46 118
rect 50 120 56 122
rect 50 118 52 120
rect 54 118 56 120
rect 50 116 56 118
rect 40 111 42 116
rect 53 111 55 116
rect 60 111 62 124
rect 80 111 82 124
rect 90 122 92 133
rect 100 122 102 126
rect 86 120 92 122
rect 86 118 88 120
rect 90 118 92 120
rect 86 116 92 118
rect 96 120 102 122
rect 96 118 98 120
rect 100 118 102 120
rect 96 116 102 118
rect 87 111 89 116
rect 100 111 102 116
rect 120 122 122 126
rect 130 122 132 133
rect 140 130 142 133
rect 140 128 146 130
rect 140 126 142 128
rect 144 126 146 128
rect 140 124 146 126
rect 154 128 160 130
rect 154 126 156 128
rect 158 126 160 128
rect 205 153 207 157
rect 185 144 187 148
rect 195 144 197 148
rect 293 153 295 157
rect 244 144 246 148
rect 254 146 256 151
rect 264 146 266 151
rect 154 124 160 126
rect 120 120 126 122
rect 120 118 122 120
rect 124 118 126 120
rect 120 116 126 118
rect 130 120 136 122
rect 130 118 132 120
rect 134 118 136 120
rect 130 116 136 118
rect 120 111 122 116
rect 133 111 135 116
rect 140 111 142 124
rect 158 123 160 124
rect 169 123 171 126
rect 185 123 187 126
rect 158 121 171 123
rect 177 121 187 123
rect 195 122 197 126
rect 205 123 207 126
rect 161 113 163 121
rect 177 117 179 121
rect 170 115 179 117
rect 191 120 197 122
rect 191 118 193 120
rect 195 118 197 120
rect 191 116 197 118
rect 201 121 207 123
rect 201 119 203 121
rect 205 119 207 121
rect 201 117 207 119
rect 244 122 246 126
rect 254 122 256 133
rect 264 130 266 133
rect 264 128 270 130
rect 264 126 266 128
rect 268 126 270 128
rect 264 124 270 126
rect 278 128 284 130
rect 278 126 280 128
rect 282 126 284 128
rect 329 153 331 157
rect 309 144 311 148
rect 319 144 321 148
rect 370 145 372 150
rect 380 145 382 150
rect 457 152 459 156
rect 390 143 392 147
rect 410 145 412 150
rect 420 145 422 150
rect 370 129 372 132
rect 366 127 372 129
rect 278 124 284 126
rect 244 120 250 122
rect 244 118 246 120
rect 248 118 250 120
rect 170 113 172 115
rect 174 113 179 115
rect 40 98 42 102
rect 53 95 55 100
rect 60 95 62 100
rect 80 95 82 100
rect 87 95 89 100
rect 100 98 102 102
rect 120 98 122 102
rect 170 111 179 113
rect 195 113 197 116
rect 177 108 179 111
rect 187 108 189 112
rect 195 111 199 113
rect 197 108 199 111
rect 204 108 206 117
rect 244 116 250 118
rect 254 120 260 122
rect 254 118 256 120
rect 258 118 260 120
rect 254 116 260 118
rect 244 111 246 116
rect 257 111 259 116
rect 264 111 266 124
rect 282 123 284 124
rect 293 123 295 126
rect 309 123 311 126
rect 282 121 295 123
rect 301 121 311 123
rect 319 122 321 126
rect 329 123 331 126
rect 366 125 368 127
rect 370 125 372 127
rect 366 123 372 125
rect 285 113 287 121
rect 301 117 303 121
rect 294 115 303 117
rect 315 120 321 122
rect 315 118 317 120
rect 319 118 321 120
rect 315 116 321 118
rect 325 121 331 123
rect 325 119 327 121
rect 329 119 331 121
rect 325 117 331 119
rect 294 113 296 115
rect 298 113 303 115
rect 161 101 163 104
rect 133 95 135 100
rect 140 95 142 100
rect 161 99 166 101
rect 164 91 166 99
rect 177 95 179 99
rect 187 91 189 99
rect 244 98 246 102
rect 294 111 303 113
rect 319 113 321 116
rect 301 108 303 111
rect 311 108 313 112
rect 319 111 323 113
rect 321 108 323 111
rect 328 108 330 117
rect 370 110 372 123
rect 380 121 382 132
rect 430 143 432 147
rect 410 129 412 132
rect 406 127 412 129
rect 406 125 408 127
rect 410 125 412 127
rect 390 121 392 125
rect 406 123 412 125
rect 376 119 382 121
rect 376 117 378 119
rect 380 117 382 119
rect 376 115 382 117
rect 386 119 392 121
rect 386 117 388 119
rect 390 117 392 119
rect 386 115 392 117
rect 377 110 379 115
rect 390 110 392 115
rect 410 110 412 123
rect 420 121 422 132
rect 493 152 495 156
rect 467 143 469 147
rect 477 143 479 147
rect 522 145 524 150
rect 532 145 534 150
rect 542 143 544 147
rect 575 145 577 150
rect 585 145 587 150
rect 662 152 664 156
rect 522 129 524 132
rect 504 127 510 129
rect 504 125 506 127
rect 508 125 510 127
rect 430 121 432 125
rect 416 119 422 121
rect 416 117 418 119
rect 420 117 422 119
rect 416 115 422 117
rect 426 119 432 121
rect 426 117 428 119
rect 430 117 432 119
rect 426 115 432 117
rect 457 122 459 125
rect 457 120 463 122
rect 457 118 459 120
rect 461 118 463 120
rect 457 116 463 118
rect 467 121 469 125
rect 477 122 479 125
rect 493 122 495 125
rect 504 123 510 125
rect 518 127 524 129
rect 518 125 520 127
rect 522 125 524 127
rect 518 123 524 125
rect 504 122 506 123
rect 467 119 473 121
rect 477 120 487 122
rect 493 120 506 122
rect 467 117 469 119
rect 471 117 473 119
rect 417 110 419 115
rect 430 110 432 115
rect 285 101 287 104
rect 197 91 199 96
rect 204 91 206 96
rect 164 89 189 91
rect 257 95 259 100
rect 264 95 266 100
rect 285 99 290 101
rect 288 91 290 99
rect 301 95 303 99
rect 311 91 313 99
rect 321 91 323 96
rect 328 91 330 96
rect 370 94 372 99
rect 377 94 379 99
rect 288 89 313 91
rect 390 97 392 101
rect 458 107 460 116
rect 467 115 473 117
rect 485 116 487 120
rect 467 112 469 115
rect 465 110 469 112
rect 485 114 494 116
rect 485 112 490 114
rect 492 112 494 114
rect 501 112 503 120
rect 465 107 467 110
rect 475 107 477 111
rect 485 110 494 112
rect 485 107 487 110
rect 410 94 412 99
rect 417 94 419 99
rect 430 97 432 101
rect 522 110 524 123
rect 532 121 534 132
rect 595 143 597 147
rect 615 145 617 150
rect 625 145 627 150
rect 575 129 577 132
rect 571 127 577 129
rect 571 125 573 127
rect 575 125 577 127
rect 542 121 544 125
rect 571 123 577 125
rect 528 119 534 121
rect 528 117 530 119
rect 532 117 534 119
rect 528 115 534 117
rect 538 119 544 121
rect 538 117 540 119
rect 542 117 544 119
rect 538 115 544 117
rect 529 110 531 115
rect 542 110 544 115
rect 575 110 577 123
rect 585 121 587 132
rect 635 143 637 147
rect 615 129 617 132
rect 611 127 617 129
rect 611 125 613 127
rect 615 125 617 127
rect 595 121 597 125
rect 611 123 617 125
rect 581 119 587 121
rect 581 117 583 119
rect 585 117 587 119
rect 581 115 587 117
rect 591 119 597 121
rect 591 117 593 119
rect 595 117 597 119
rect 591 115 597 117
rect 582 110 584 115
rect 595 110 597 115
rect 615 110 617 123
rect 625 121 627 132
rect 698 152 700 156
rect 672 143 674 147
rect 682 143 684 147
rect 727 145 729 150
rect 737 145 739 150
rect 795 153 797 157
rect 802 153 804 157
rect 747 143 749 147
rect 782 143 784 148
rect 727 129 729 132
rect 709 127 715 129
rect 709 125 711 127
rect 713 125 715 127
rect 635 121 637 125
rect 621 119 627 121
rect 621 117 623 119
rect 625 117 627 119
rect 621 115 627 117
rect 631 119 637 121
rect 631 117 633 119
rect 635 117 637 119
rect 631 115 637 117
rect 662 122 664 125
rect 662 120 668 122
rect 662 118 664 120
rect 666 118 668 120
rect 662 116 668 118
rect 672 121 674 125
rect 682 122 684 125
rect 698 122 700 125
rect 709 123 715 125
rect 723 127 729 129
rect 723 125 725 127
rect 727 125 729 127
rect 723 123 729 125
rect 709 122 711 123
rect 672 119 678 121
rect 682 120 692 122
rect 698 120 711 122
rect 672 117 674 119
rect 676 117 678 119
rect 622 110 624 115
rect 635 110 637 115
rect 501 100 503 103
rect 498 98 503 100
rect 458 90 460 95
rect 465 90 467 95
rect 475 90 477 98
rect 485 94 487 98
rect 498 90 500 98
rect 475 88 500 90
rect 522 94 524 99
rect 529 94 531 99
rect 542 97 544 101
rect 575 94 577 99
rect 582 94 584 99
rect 595 97 597 101
rect 663 107 665 116
rect 672 115 678 117
rect 690 116 692 120
rect 672 112 674 115
rect 670 110 674 112
rect 690 114 699 116
rect 690 112 695 114
rect 697 112 699 114
rect 706 112 708 120
rect 670 107 672 110
rect 680 107 682 111
rect 690 110 699 112
rect 690 107 692 110
rect 615 94 617 99
rect 622 94 624 99
rect 635 97 637 101
rect 727 110 729 123
rect 737 121 739 132
rect 871 153 873 157
rect 822 144 824 148
rect 832 146 834 151
rect 842 146 844 151
rect 747 121 749 125
rect 733 119 739 121
rect 733 117 735 119
rect 737 117 739 119
rect 733 115 739 117
rect 743 119 749 121
rect 743 117 745 119
rect 747 117 749 119
rect 743 115 749 117
rect 734 110 736 115
rect 747 110 749 115
rect 782 122 784 125
rect 795 122 797 132
rect 802 129 804 132
rect 802 127 808 129
rect 802 125 804 127
rect 806 125 808 127
rect 802 123 808 125
rect 782 120 788 122
rect 782 118 784 120
rect 786 118 788 120
rect 782 116 788 118
rect 792 120 798 122
rect 792 118 794 120
rect 796 118 798 120
rect 792 116 798 118
rect 782 113 784 116
rect 792 113 794 116
rect 802 113 804 123
rect 822 122 824 126
rect 832 122 834 133
rect 842 130 844 133
rect 842 128 848 130
rect 842 126 844 128
rect 846 126 848 128
rect 842 124 848 126
rect 856 128 862 130
rect 856 126 858 128
rect 860 126 862 128
rect 907 153 909 157
rect 887 144 889 148
rect 897 144 899 148
rect 976 153 978 157
rect 927 144 929 148
rect 937 146 939 151
rect 947 146 949 151
rect 856 124 862 126
rect 822 120 828 122
rect 822 118 824 120
rect 826 118 828 120
rect 822 116 828 118
rect 832 120 838 122
rect 832 118 834 120
rect 836 118 838 120
rect 832 116 838 118
rect 706 100 708 103
rect 703 98 708 100
rect 822 111 824 116
rect 835 111 837 116
rect 842 111 844 124
rect 860 123 862 124
rect 871 123 873 126
rect 887 123 889 126
rect 860 121 873 123
rect 879 121 889 123
rect 897 122 899 126
rect 907 123 909 126
rect 863 113 865 121
rect 879 117 881 121
rect 872 115 881 117
rect 893 120 899 122
rect 893 118 895 120
rect 897 118 899 120
rect 893 116 899 118
rect 903 121 909 123
rect 903 119 905 121
rect 907 119 909 121
rect 903 117 909 119
rect 927 122 929 126
rect 937 122 939 133
rect 947 130 949 133
rect 947 128 953 130
rect 947 126 949 128
rect 951 126 953 128
rect 947 124 953 126
rect 961 128 967 130
rect 961 126 963 128
rect 965 126 967 128
rect 1012 153 1014 157
rect 992 144 994 148
rect 1002 144 1004 148
rect 1045 153 1047 157
rect 1052 153 1054 157
rect 1032 143 1034 148
rect 961 124 967 126
rect 927 120 933 122
rect 927 118 929 120
rect 931 118 933 120
rect 872 113 874 115
rect 876 113 881 115
rect 663 90 665 95
rect 670 90 672 95
rect 680 90 682 98
rect 690 94 692 98
rect 703 90 705 98
rect 680 88 705 90
rect 727 94 729 99
rect 734 94 736 99
rect 747 97 749 101
rect 782 99 784 104
rect 792 102 794 107
rect 802 102 804 107
rect 822 98 824 102
rect 872 111 881 113
rect 897 113 899 116
rect 879 108 881 111
rect 889 108 891 112
rect 897 111 901 113
rect 899 108 901 111
rect 906 108 908 117
rect 927 116 933 118
rect 937 120 943 122
rect 937 118 939 120
rect 941 118 943 120
rect 937 116 943 118
rect 927 111 929 116
rect 940 111 942 116
rect 947 111 949 124
rect 965 123 967 124
rect 976 123 978 126
rect 992 123 994 126
rect 965 121 978 123
rect 984 121 994 123
rect 1002 122 1004 126
rect 1012 123 1014 126
rect 1121 153 1123 157
rect 1072 144 1074 148
rect 1082 146 1084 151
rect 1092 146 1094 151
rect 968 113 970 121
rect 984 117 986 121
rect 977 115 986 117
rect 998 120 1004 122
rect 998 118 1000 120
rect 1002 118 1004 120
rect 998 116 1004 118
rect 1008 121 1014 123
rect 1008 119 1010 121
rect 1012 119 1014 121
rect 1008 117 1014 119
rect 1032 122 1034 125
rect 1045 122 1047 132
rect 1052 129 1054 132
rect 1052 127 1058 129
rect 1052 125 1054 127
rect 1056 125 1058 127
rect 1052 123 1058 125
rect 1032 120 1038 122
rect 1032 118 1034 120
rect 1036 118 1038 120
rect 977 113 979 115
rect 981 113 986 115
rect 863 101 865 104
rect 835 95 837 100
rect 842 95 844 100
rect 863 99 868 101
rect 866 91 868 99
rect 879 95 881 99
rect 889 91 891 99
rect 927 98 929 102
rect 977 111 986 113
rect 1002 113 1004 116
rect 984 108 986 111
rect 994 108 996 112
rect 1002 111 1006 113
rect 1004 108 1006 111
rect 1011 108 1013 117
rect 1032 116 1038 118
rect 1042 120 1048 122
rect 1042 118 1044 120
rect 1046 118 1048 120
rect 1042 116 1048 118
rect 1032 113 1034 116
rect 1042 113 1044 116
rect 1052 113 1054 123
rect 1072 122 1074 126
rect 1082 122 1084 133
rect 1092 130 1094 133
rect 1092 128 1098 130
rect 1092 126 1094 128
rect 1096 126 1098 128
rect 1092 124 1098 126
rect 1106 128 1112 130
rect 1106 126 1108 128
rect 1110 126 1112 128
rect 1157 153 1159 157
rect 1137 144 1139 148
rect 1147 144 1149 148
rect 1226 153 1228 157
rect 1177 144 1179 148
rect 1187 146 1189 151
rect 1197 146 1199 151
rect 1106 124 1112 126
rect 1072 120 1078 122
rect 1072 118 1074 120
rect 1076 118 1078 120
rect 1072 116 1078 118
rect 1082 120 1088 122
rect 1082 118 1084 120
rect 1086 118 1088 120
rect 1082 116 1088 118
rect 968 101 970 104
rect 899 91 901 96
rect 906 91 908 96
rect 866 89 891 91
rect 940 95 942 100
rect 947 95 949 100
rect 968 99 973 101
rect 971 91 973 99
rect 984 95 986 99
rect 994 91 996 99
rect 1072 111 1074 116
rect 1085 111 1087 116
rect 1092 111 1094 124
rect 1110 123 1112 124
rect 1121 123 1123 126
rect 1137 123 1139 126
rect 1110 121 1123 123
rect 1129 121 1139 123
rect 1147 122 1149 126
rect 1157 123 1159 126
rect 1113 113 1115 121
rect 1129 117 1131 121
rect 1122 115 1131 117
rect 1143 120 1149 122
rect 1143 118 1145 120
rect 1147 118 1149 120
rect 1143 116 1149 118
rect 1153 121 1159 123
rect 1153 119 1155 121
rect 1157 119 1159 121
rect 1153 117 1159 119
rect 1177 122 1179 126
rect 1187 122 1189 133
rect 1197 130 1199 133
rect 1197 128 1203 130
rect 1197 126 1199 128
rect 1201 126 1203 128
rect 1197 124 1203 126
rect 1211 128 1217 130
rect 1211 126 1213 128
rect 1215 126 1217 128
rect 1262 153 1264 157
rect 1242 144 1244 148
rect 1252 144 1254 148
rect 1295 153 1297 157
rect 1302 153 1304 157
rect 1282 143 1284 148
rect 1211 124 1217 126
rect 1177 120 1183 122
rect 1177 118 1179 120
rect 1181 118 1183 120
rect 1122 113 1124 115
rect 1126 113 1131 115
rect 1032 99 1034 104
rect 1042 102 1044 107
rect 1052 102 1054 107
rect 1004 91 1006 96
rect 1011 91 1013 96
rect 971 89 996 91
rect 1072 98 1074 102
rect 1122 111 1131 113
rect 1147 113 1149 116
rect 1129 108 1131 111
rect 1139 108 1141 112
rect 1147 111 1151 113
rect 1149 108 1151 111
rect 1156 108 1158 117
rect 1177 116 1183 118
rect 1187 120 1193 122
rect 1187 118 1189 120
rect 1191 118 1193 120
rect 1187 116 1193 118
rect 1177 111 1179 116
rect 1190 111 1192 116
rect 1197 111 1199 124
rect 1215 123 1217 124
rect 1226 123 1228 126
rect 1242 123 1244 126
rect 1215 121 1228 123
rect 1234 121 1244 123
rect 1252 122 1254 126
rect 1262 123 1264 126
rect 1371 153 1373 157
rect 1322 144 1324 148
rect 1332 146 1334 151
rect 1342 146 1344 151
rect 1218 113 1220 121
rect 1234 117 1236 121
rect 1227 115 1236 117
rect 1248 120 1254 122
rect 1248 118 1250 120
rect 1252 118 1254 120
rect 1248 116 1254 118
rect 1258 121 1264 123
rect 1258 119 1260 121
rect 1262 119 1264 121
rect 1258 117 1264 119
rect 1282 122 1284 125
rect 1295 122 1297 132
rect 1302 129 1304 132
rect 1302 127 1308 129
rect 1302 125 1304 127
rect 1306 125 1308 127
rect 1302 123 1308 125
rect 1282 120 1288 122
rect 1282 118 1284 120
rect 1286 118 1288 120
rect 1227 113 1229 115
rect 1231 113 1236 115
rect 1113 101 1115 104
rect 1085 95 1087 100
rect 1092 95 1094 100
rect 1113 99 1118 101
rect 1116 91 1118 99
rect 1129 95 1131 99
rect 1139 91 1141 99
rect 1177 98 1179 102
rect 1227 111 1236 113
rect 1252 113 1254 116
rect 1234 108 1236 111
rect 1244 108 1246 112
rect 1252 111 1256 113
rect 1254 108 1256 111
rect 1261 108 1263 117
rect 1282 116 1288 118
rect 1292 120 1298 122
rect 1292 118 1294 120
rect 1296 118 1298 120
rect 1292 116 1298 118
rect 1282 113 1284 116
rect 1292 113 1294 116
rect 1302 113 1304 123
rect 1322 122 1324 126
rect 1332 122 1334 133
rect 1342 130 1344 133
rect 1342 128 1348 130
rect 1342 126 1344 128
rect 1346 126 1348 128
rect 1342 124 1348 126
rect 1356 128 1362 130
rect 1356 126 1358 128
rect 1360 126 1362 128
rect 1407 153 1409 157
rect 1387 144 1389 148
rect 1397 144 1399 148
rect 1476 153 1478 157
rect 1427 144 1429 148
rect 1437 146 1439 151
rect 1447 146 1449 151
rect 1356 124 1362 126
rect 1322 120 1328 122
rect 1322 118 1324 120
rect 1326 118 1328 120
rect 1322 116 1328 118
rect 1332 120 1338 122
rect 1332 118 1334 120
rect 1336 118 1338 120
rect 1332 116 1338 118
rect 1218 101 1220 104
rect 1149 91 1151 96
rect 1156 91 1158 96
rect 1116 89 1141 91
rect 1190 95 1192 100
rect 1197 95 1199 100
rect 1218 99 1223 101
rect 1221 91 1223 99
rect 1234 95 1236 99
rect 1244 91 1246 99
rect 1322 111 1324 116
rect 1335 111 1337 116
rect 1342 111 1344 124
rect 1360 123 1362 124
rect 1371 123 1373 126
rect 1387 123 1389 126
rect 1360 121 1373 123
rect 1379 121 1389 123
rect 1397 122 1399 126
rect 1407 123 1409 126
rect 1363 113 1365 121
rect 1379 117 1381 121
rect 1372 115 1381 117
rect 1393 120 1399 122
rect 1393 118 1395 120
rect 1397 118 1399 120
rect 1393 116 1399 118
rect 1403 121 1409 123
rect 1403 119 1405 121
rect 1407 119 1409 121
rect 1403 117 1409 119
rect 1427 122 1429 126
rect 1437 122 1439 133
rect 1447 130 1449 133
rect 1447 128 1453 130
rect 1447 126 1449 128
rect 1451 126 1453 128
rect 1447 124 1453 126
rect 1461 128 1467 130
rect 1461 126 1463 128
rect 1465 126 1467 128
rect 1512 153 1514 157
rect 1492 144 1494 148
rect 1502 144 1504 148
rect 1545 153 1547 157
rect 1552 153 1554 157
rect 1532 143 1534 148
rect 1461 124 1467 126
rect 1427 120 1433 122
rect 1427 118 1429 120
rect 1431 118 1433 120
rect 1372 113 1374 115
rect 1376 113 1381 115
rect 1282 99 1284 104
rect 1292 102 1294 107
rect 1302 102 1304 107
rect 1254 91 1256 96
rect 1261 91 1263 96
rect 1221 89 1246 91
rect 1322 98 1324 102
rect 1372 111 1381 113
rect 1397 113 1399 116
rect 1379 108 1381 111
rect 1389 108 1391 112
rect 1397 111 1401 113
rect 1399 108 1401 111
rect 1406 108 1408 117
rect 1427 116 1433 118
rect 1437 120 1443 122
rect 1437 118 1439 120
rect 1441 118 1443 120
rect 1437 116 1443 118
rect 1427 111 1429 116
rect 1440 111 1442 116
rect 1447 111 1449 124
rect 1465 123 1467 124
rect 1476 123 1478 126
rect 1492 123 1494 126
rect 1465 121 1478 123
rect 1484 121 1494 123
rect 1502 122 1504 126
rect 1512 123 1514 126
rect 1621 153 1623 157
rect 1572 144 1574 148
rect 1582 146 1584 151
rect 1592 146 1594 151
rect 1468 113 1470 121
rect 1484 117 1486 121
rect 1477 115 1486 117
rect 1498 120 1504 122
rect 1498 118 1500 120
rect 1502 118 1504 120
rect 1498 116 1504 118
rect 1508 121 1514 123
rect 1508 119 1510 121
rect 1512 119 1514 121
rect 1508 117 1514 119
rect 1532 122 1534 125
rect 1545 122 1547 132
rect 1552 129 1554 132
rect 1552 127 1558 129
rect 1552 125 1554 127
rect 1556 125 1558 127
rect 1552 123 1558 125
rect 1532 120 1538 122
rect 1532 118 1534 120
rect 1536 118 1538 120
rect 1477 113 1479 115
rect 1481 113 1486 115
rect 1363 101 1365 104
rect 1335 95 1337 100
rect 1342 95 1344 100
rect 1363 99 1368 101
rect 1366 91 1368 99
rect 1379 95 1381 99
rect 1389 91 1391 99
rect 1427 98 1429 102
rect 1477 111 1486 113
rect 1502 113 1504 116
rect 1484 108 1486 111
rect 1494 108 1496 112
rect 1502 111 1506 113
rect 1504 108 1506 111
rect 1511 108 1513 117
rect 1532 116 1538 118
rect 1542 120 1548 122
rect 1542 118 1544 120
rect 1546 118 1548 120
rect 1542 116 1548 118
rect 1532 113 1534 116
rect 1542 113 1544 116
rect 1552 113 1554 123
rect 1572 122 1574 126
rect 1582 122 1584 133
rect 1592 130 1594 133
rect 1592 128 1598 130
rect 1592 126 1594 128
rect 1596 126 1598 128
rect 1592 124 1598 126
rect 1606 128 1612 130
rect 1606 126 1608 128
rect 1610 126 1612 128
rect 1657 153 1659 157
rect 1637 144 1639 148
rect 1647 144 1649 148
rect 1726 153 1728 157
rect 1677 144 1679 148
rect 1687 146 1689 151
rect 1697 146 1699 151
rect 1606 124 1612 126
rect 1572 120 1578 122
rect 1572 118 1574 120
rect 1576 118 1578 120
rect 1572 116 1578 118
rect 1582 120 1588 122
rect 1582 118 1584 120
rect 1586 118 1588 120
rect 1582 116 1588 118
rect 1468 101 1470 104
rect 1399 91 1401 96
rect 1406 91 1408 96
rect 1366 89 1391 91
rect 1440 95 1442 100
rect 1447 95 1449 100
rect 1468 99 1473 101
rect 1471 91 1473 99
rect 1484 95 1486 99
rect 1494 91 1496 99
rect 1572 111 1574 116
rect 1585 111 1587 116
rect 1592 111 1594 124
rect 1610 123 1612 124
rect 1621 123 1623 126
rect 1637 123 1639 126
rect 1610 121 1623 123
rect 1629 121 1639 123
rect 1647 122 1649 126
rect 1657 123 1659 126
rect 1613 113 1615 121
rect 1629 117 1631 121
rect 1622 115 1631 117
rect 1643 120 1649 122
rect 1643 118 1645 120
rect 1647 118 1649 120
rect 1643 116 1649 118
rect 1653 121 1659 123
rect 1653 119 1655 121
rect 1657 119 1659 121
rect 1653 117 1659 119
rect 1677 122 1679 126
rect 1687 122 1689 133
rect 1697 130 1699 133
rect 1697 128 1703 130
rect 1697 126 1699 128
rect 1701 126 1703 128
rect 1697 124 1703 126
rect 1711 128 1717 130
rect 1711 126 1713 128
rect 1715 126 1717 128
rect 1762 153 1764 157
rect 1742 144 1744 148
rect 1752 144 1754 148
rect 1830 144 1832 148
rect 1840 146 1842 151
rect 1850 146 1852 151
rect 1870 146 1872 151
rect 1880 146 1882 151
rect 1959 153 1961 157
rect 1890 144 1892 148
rect 1910 144 1912 148
rect 1920 146 1922 151
rect 1930 146 1932 151
rect 1711 124 1717 126
rect 1677 120 1683 122
rect 1677 118 1679 120
rect 1681 118 1683 120
rect 1622 113 1624 115
rect 1626 113 1631 115
rect 1532 99 1534 104
rect 1542 102 1544 107
rect 1552 102 1554 107
rect 1504 91 1506 96
rect 1511 91 1513 96
rect 1471 89 1496 91
rect 1572 98 1574 102
rect 1622 111 1631 113
rect 1647 113 1649 116
rect 1629 108 1631 111
rect 1639 108 1641 112
rect 1647 111 1651 113
rect 1649 108 1651 111
rect 1656 108 1658 117
rect 1677 116 1683 118
rect 1687 120 1693 122
rect 1687 118 1689 120
rect 1691 118 1693 120
rect 1687 116 1693 118
rect 1677 111 1679 116
rect 1690 111 1692 116
rect 1697 111 1699 124
rect 1715 123 1717 124
rect 1726 123 1728 126
rect 1742 123 1744 126
rect 1715 121 1728 123
rect 1734 121 1744 123
rect 1752 122 1754 126
rect 1762 123 1764 126
rect 1718 113 1720 121
rect 1734 117 1736 121
rect 1727 115 1736 117
rect 1748 120 1754 122
rect 1748 118 1750 120
rect 1752 118 1754 120
rect 1748 116 1754 118
rect 1758 121 1764 123
rect 1758 119 1760 121
rect 1762 119 1764 121
rect 1758 117 1764 119
rect 1830 122 1832 126
rect 1840 122 1842 133
rect 1850 130 1852 133
rect 1870 130 1872 133
rect 1850 128 1856 130
rect 1850 126 1852 128
rect 1854 126 1856 128
rect 1850 124 1856 126
rect 1866 128 1872 130
rect 1866 126 1868 128
rect 1870 126 1872 128
rect 1866 124 1872 126
rect 1830 120 1836 122
rect 1830 118 1832 120
rect 1834 118 1836 120
rect 1727 113 1729 115
rect 1731 113 1736 115
rect 1613 101 1615 104
rect 1585 95 1587 100
rect 1592 95 1594 100
rect 1613 99 1618 101
rect 1616 91 1618 99
rect 1629 95 1631 99
rect 1639 91 1641 99
rect 1677 98 1679 102
rect 1727 111 1736 113
rect 1752 113 1754 116
rect 1734 108 1736 111
rect 1744 108 1746 112
rect 1752 111 1756 113
rect 1754 108 1756 111
rect 1761 108 1763 117
rect 1830 116 1836 118
rect 1840 120 1846 122
rect 1840 118 1842 120
rect 1844 118 1846 120
rect 1840 116 1846 118
rect 1830 111 1832 116
rect 1843 111 1845 116
rect 1850 111 1852 124
rect 1870 111 1872 124
rect 1880 122 1882 133
rect 1890 122 1892 126
rect 1876 120 1882 122
rect 1876 118 1878 120
rect 1880 118 1882 120
rect 1876 116 1882 118
rect 1886 120 1892 122
rect 1886 118 1888 120
rect 1890 118 1892 120
rect 1886 116 1892 118
rect 1877 111 1879 116
rect 1890 111 1892 116
rect 1910 122 1912 126
rect 1920 122 1922 133
rect 1930 130 1932 133
rect 1930 128 1936 130
rect 1930 126 1932 128
rect 1934 126 1936 128
rect 1930 124 1936 126
rect 1944 128 1950 130
rect 1944 126 1946 128
rect 1948 126 1950 128
rect 1995 153 1997 157
rect 1975 144 1977 148
rect 1985 144 1987 148
rect 1944 124 1950 126
rect 1910 120 1916 122
rect 1910 118 1912 120
rect 1914 118 1916 120
rect 1910 116 1916 118
rect 1920 120 1926 122
rect 1920 118 1922 120
rect 1924 118 1926 120
rect 1920 116 1926 118
rect 1910 111 1912 116
rect 1923 111 1925 116
rect 1930 111 1932 124
rect 1948 123 1950 124
rect 1959 123 1961 126
rect 1975 123 1977 126
rect 1948 121 1961 123
rect 1967 121 1977 123
rect 1985 122 1987 126
rect 1995 123 1997 126
rect 1951 113 1953 121
rect 1967 117 1969 121
rect 1960 115 1969 117
rect 1981 120 1987 122
rect 1981 118 1983 120
rect 1985 118 1987 120
rect 1981 116 1987 118
rect 1991 121 1997 123
rect 1991 119 1993 121
rect 1995 119 1997 121
rect 1991 117 1997 119
rect 1960 113 1962 115
rect 1964 113 1969 115
rect 1718 101 1720 104
rect 1649 91 1651 96
rect 1656 91 1658 96
rect 1616 89 1641 91
rect 1690 95 1692 100
rect 1697 95 1699 100
rect 1718 99 1723 101
rect 1721 91 1723 99
rect 1734 95 1736 99
rect 1744 91 1746 99
rect 1830 98 1832 102
rect 1754 91 1756 96
rect 1761 91 1763 96
rect 1721 89 1746 91
rect 1843 95 1845 100
rect 1850 95 1852 100
rect 1870 95 1872 100
rect 1877 95 1879 100
rect 1890 98 1892 102
rect 1910 98 1912 102
rect 1960 111 1969 113
rect 1985 113 1987 116
rect 1967 108 1969 111
rect 1977 108 1979 112
rect 1985 111 1989 113
rect 1987 108 1989 111
rect 1994 108 1996 117
rect 1951 101 1953 104
rect 1923 95 1925 100
rect 1930 95 1932 100
rect 1951 99 1956 101
rect 1954 91 1956 99
rect 1967 95 1969 99
rect 1977 91 1979 99
rect 1987 91 1989 96
rect 1994 91 1996 96
rect 1954 89 1979 91
rect 14 60 16 65
rect 24 57 26 62
rect 34 57 36 62
rect 54 62 56 66
rect 67 64 69 69
rect 74 64 76 69
rect 98 73 123 75
rect 98 65 100 73
rect 111 65 113 69
rect 121 65 123 73
rect 131 68 133 73
rect 138 68 140 73
rect 95 63 100 65
rect 95 60 97 63
rect 14 48 16 51
rect 24 48 26 51
rect 14 46 20 48
rect 14 44 16 46
rect 18 44 20 46
rect 14 42 20 44
rect 24 46 30 48
rect 24 44 26 46
rect 28 44 30 46
rect 24 42 30 44
rect 14 39 16 42
rect 27 32 29 42
rect 34 41 36 51
rect 54 48 56 53
rect 67 48 69 53
rect 54 46 60 48
rect 54 44 56 46
rect 58 44 60 46
rect 54 42 60 44
rect 64 46 70 48
rect 64 44 66 46
rect 68 44 70 46
rect 64 42 70 44
rect 34 39 40 41
rect 34 37 36 39
rect 38 37 40 39
rect 54 38 56 42
rect 34 35 40 37
rect 34 32 36 35
rect 14 16 16 21
rect 64 31 66 42
rect 74 40 76 53
rect 159 62 161 66
rect 172 64 174 69
rect 179 64 181 69
rect 203 73 228 75
rect 203 65 205 73
rect 216 65 218 69
rect 226 65 228 73
rect 236 68 238 73
rect 243 68 245 73
rect 111 53 113 56
rect 104 51 113 53
rect 121 52 123 56
rect 131 53 133 56
rect 95 43 97 51
rect 104 49 106 51
rect 108 49 113 51
rect 104 47 113 49
rect 129 51 133 53
rect 129 48 131 51
rect 111 43 113 47
rect 125 46 131 48
rect 138 47 140 56
rect 200 63 205 65
rect 200 60 202 63
rect 159 48 161 53
rect 172 48 174 53
rect 125 44 127 46
rect 129 44 131 46
rect 92 41 105 43
rect 111 41 121 43
rect 125 42 131 44
rect 92 40 94 41
rect 74 38 80 40
rect 74 36 76 38
rect 78 36 80 38
rect 74 34 80 36
rect 88 38 94 40
rect 103 38 105 41
rect 119 38 121 41
rect 129 38 131 42
rect 135 45 141 47
rect 135 43 137 45
rect 139 43 141 45
rect 135 41 141 43
rect 139 38 141 41
rect 159 46 165 48
rect 159 44 161 46
rect 163 44 165 46
rect 159 42 165 44
rect 169 46 175 48
rect 169 44 171 46
rect 173 44 175 46
rect 169 42 175 44
rect 159 38 161 42
rect 88 36 90 38
rect 92 36 94 38
rect 88 34 94 36
rect 74 31 76 34
rect 54 16 56 20
rect 64 13 66 18
rect 74 13 76 18
rect 27 7 29 11
rect 34 7 36 11
rect 119 16 121 20
rect 129 16 131 20
rect 103 7 105 11
rect 169 31 171 42
rect 179 40 181 53
rect 264 60 266 65
rect 216 53 218 56
rect 209 51 218 53
rect 226 52 228 56
rect 236 53 238 56
rect 200 43 202 51
rect 209 49 211 51
rect 213 49 218 51
rect 209 47 218 49
rect 234 51 238 53
rect 234 48 236 51
rect 216 43 218 47
rect 230 46 236 48
rect 243 47 245 56
rect 274 57 276 62
rect 284 57 286 62
rect 304 62 306 66
rect 317 64 319 69
rect 324 64 326 69
rect 348 73 373 75
rect 348 65 350 73
rect 361 65 363 69
rect 371 65 373 73
rect 381 68 383 73
rect 388 68 390 73
rect 345 63 350 65
rect 345 60 347 63
rect 264 48 266 51
rect 274 48 276 51
rect 230 44 232 46
rect 234 44 236 46
rect 197 41 210 43
rect 216 41 226 43
rect 230 42 236 44
rect 197 40 199 41
rect 179 38 185 40
rect 179 36 181 38
rect 183 36 185 38
rect 179 34 185 36
rect 193 38 199 40
rect 208 38 210 41
rect 224 38 226 41
rect 234 38 236 42
rect 240 45 246 47
rect 240 43 242 45
rect 244 43 246 45
rect 240 41 246 43
rect 244 38 246 41
rect 264 46 270 48
rect 264 44 266 46
rect 268 44 270 46
rect 264 42 270 44
rect 274 46 280 48
rect 274 44 276 46
rect 278 44 280 46
rect 274 42 280 44
rect 264 39 266 42
rect 193 36 195 38
rect 197 36 199 38
rect 193 34 199 36
rect 179 31 181 34
rect 159 16 161 20
rect 169 13 171 18
rect 179 13 181 18
rect 139 7 141 11
rect 224 16 226 20
rect 234 16 236 20
rect 208 7 210 11
rect 277 32 279 42
rect 284 41 286 51
rect 304 48 306 53
rect 317 48 319 53
rect 304 46 310 48
rect 304 44 306 46
rect 308 44 310 46
rect 304 42 310 44
rect 314 46 320 48
rect 314 44 316 46
rect 318 44 320 46
rect 314 42 320 44
rect 284 39 290 41
rect 284 37 286 39
rect 288 37 290 39
rect 304 38 306 42
rect 284 35 290 37
rect 284 32 286 35
rect 264 16 266 21
rect 244 7 246 11
rect 314 31 316 42
rect 324 40 326 53
rect 409 62 411 66
rect 422 64 424 69
rect 429 64 431 69
rect 453 73 478 75
rect 453 65 455 73
rect 466 65 468 69
rect 476 65 478 73
rect 486 68 488 73
rect 493 68 495 73
rect 361 53 363 56
rect 354 51 363 53
rect 371 52 373 56
rect 381 53 383 56
rect 345 43 347 51
rect 354 49 356 51
rect 358 49 363 51
rect 354 47 363 49
rect 379 51 383 53
rect 379 48 381 51
rect 361 43 363 47
rect 375 46 381 48
rect 388 47 390 56
rect 450 63 455 65
rect 450 60 452 63
rect 409 48 411 53
rect 422 48 424 53
rect 375 44 377 46
rect 379 44 381 46
rect 342 41 355 43
rect 361 41 371 43
rect 375 42 381 44
rect 342 40 344 41
rect 324 38 330 40
rect 324 36 326 38
rect 328 36 330 38
rect 324 34 330 36
rect 338 38 344 40
rect 353 38 355 41
rect 369 38 371 41
rect 379 38 381 42
rect 385 45 391 47
rect 385 43 387 45
rect 389 43 391 45
rect 385 41 391 43
rect 389 38 391 41
rect 409 46 415 48
rect 409 44 411 46
rect 413 44 415 46
rect 409 42 415 44
rect 419 46 425 48
rect 419 44 421 46
rect 423 44 425 46
rect 419 42 425 44
rect 409 38 411 42
rect 338 36 340 38
rect 342 36 344 38
rect 338 34 344 36
rect 324 31 326 34
rect 304 16 306 20
rect 314 13 316 18
rect 324 13 326 18
rect 277 7 279 11
rect 284 7 286 11
rect 369 16 371 20
rect 379 16 381 20
rect 353 7 355 11
rect 419 31 421 42
rect 429 40 431 53
rect 514 60 516 65
rect 466 53 468 56
rect 459 51 468 53
rect 476 52 478 56
rect 486 53 488 56
rect 450 43 452 51
rect 459 49 461 51
rect 463 49 468 51
rect 459 47 468 49
rect 484 51 488 53
rect 484 48 486 51
rect 466 43 468 47
rect 480 46 486 48
rect 493 47 495 56
rect 524 57 526 62
rect 534 57 536 62
rect 554 62 556 66
rect 567 64 569 69
rect 574 64 576 69
rect 598 73 623 75
rect 598 65 600 73
rect 611 65 613 69
rect 621 65 623 73
rect 631 68 633 73
rect 638 68 640 73
rect 595 63 600 65
rect 595 60 597 63
rect 514 48 516 51
rect 524 48 526 51
rect 480 44 482 46
rect 484 44 486 46
rect 447 41 460 43
rect 466 41 476 43
rect 480 42 486 44
rect 447 40 449 41
rect 429 38 435 40
rect 429 36 431 38
rect 433 36 435 38
rect 429 34 435 36
rect 443 38 449 40
rect 458 38 460 41
rect 474 38 476 41
rect 484 38 486 42
rect 490 45 496 47
rect 490 43 492 45
rect 494 43 496 45
rect 490 41 496 43
rect 494 38 496 41
rect 514 46 520 48
rect 514 44 516 46
rect 518 44 520 46
rect 514 42 520 44
rect 524 46 530 48
rect 524 44 526 46
rect 528 44 530 46
rect 524 42 530 44
rect 514 39 516 42
rect 443 36 445 38
rect 447 36 449 38
rect 443 34 449 36
rect 429 31 431 34
rect 409 16 411 20
rect 419 13 421 18
rect 429 13 431 18
rect 389 7 391 11
rect 474 16 476 20
rect 484 16 486 20
rect 458 7 460 11
rect 527 32 529 42
rect 534 41 536 51
rect 554 48 556 53
rect 567 48 569 53
rect 554 46 560 48
rect 554 44 556 46
rect 558 44 560 46
rect 554 42 560 44
rect 564 46 570 48
rect 564 44 566 46
rect 568 44 570 46
rect 564 42 570 44
rect 534 39 540 41
rect 534 37 536 39
rect 538 37 540 39
rect 554 38 556 42
rect 534 35 540 37
rect 534 32 536 35
rect 514 16 516 21
rect 494 7 496 11
rect 564 31 566 42
rect 574 40 576 53
rect 659 62 661 66
rect 672 64 674 69
rect 679 64 681 69
rect 703 73 728 75
rect 703 65 705 73
rect 716 65 718 69
rect 726 65 728 73
rect 736 68 738 73
rect 743 68 745 73
rect 611 53 613 56
rect 604 51 613 53
rect 621 52 623 56
rect 631 53 633 56
rect 595 43 597 51
rect 604 49 606 51
rect 608 49 613 51
rect 604 47 613 49
rect 629 51 633 53
rect 629 48 631 51
rect 611 43 613 47
rect 625 46 631 48
rect 638 47 640 56
rect 700 63 705 65
rect 700 60 702 63
rect 659 48 661 53
rect 672 48 674 53
rect 625 44 627 46
rect 629 44 631 46
rect 592 41 605 43
rect 611 41 621 43
rect 625 42 631 44
rect 592 40 594 41
rect 574 38 580 40
rect 574 36 576 38
rect 578 36 580 38
rect 574 34 580 36
rect 588 38 594 40
rect 603 38 605 41
rect 619 38 621 41
rect 629 38 631 42
rect 635 45 641 47
rect 635 43 637 45
rect 639 43 641 45
rect 635 41 641 43
rect 639 38 641 41
rect 659 46 665 48
rect 659 44 661 46
rect 663 44 665 46
rect 659 42 665 44
rect 669 46 675 48
rect 669 44 671 46
rect 673 44 675 46
rect 669 42 675 44
rect 659 38 661 42
rect 588 36 590 38
rect 592 36 594 38
rect 588 34 594 36
rect 574 31 576 34
rect 554 16 556 20
rect 564 13 566 18
rect 574 13 576 18
rect 527 7 529 11
rect 534 7 536 11
rect 619 16 621 20
rect 629 16 631 20
rect 603 7 605 11
rect 669 31 671 42
rect 679 40 681 53
rect 764 60 766 65
rect 716 53 718 56
rect 709 51 718 53
rect 726 52 728 56
rect 736 53 738 56
rect 700 43 702 51
rect 709 49 711 51
rect 713 49 718 51
rect 709 47 718 49
rect 734 51 738 53
rect 734 48 736 51
rect 716 43 718 47
rect 730 46 736 48
rect 743 47 745 56
rect 774 57 776 62
rect 784 57 786 62
rect 804 62 806 66
rect 817 64 819 69
rect 824 64 826 69
rect 848 73 873 75
rect 848 65 850 73
rect 861 65 863 69
rect 871 65 873 73
rect 881 68 883 73
rect 888 68 890 73
rect 845 63 850 65
rect 845 60 847 63
rect 764 48 766 51
rect 774 48 776 51
rect 730 44 732 46
rect 734 44 736 46
rect 697 41 710 43
rect 716 41 726 43
rect 730 42 736 44
rect 697 40 699 41
rect 679 38 685 40
rect 679 36 681 38
rect 683 36 685 38
rect 679 34 685 36
rect 693 38 699 40
rect 708 38 710 41
rect 724 38 726 41
rect 734 38 736 42
rect 740 45 746 47
rect 740 43 742 45
rect 744 43 746 45
rect 740 41 746 43
rect 744 38 746 41
rect 764 46 770 48
rect 764 44 766 46
rect 768 44 770 46
rect 764 42 770 44
rect 774 46 780 48
rect 774 44 776 46
rect 778 44 780 46
rect 774 42 780 44
rect 764 39 766 42
rect 693 36 695 38
rect 697 36 699 38
rect 693 34 699 36
rect 679 31 681 34
rect 659 16 661 20
rect 669 13 671 18
rect 679 13 681 18
rect 639 7 641 11
rect 724 16 726 20
rect 734 16 736 20
rect 708 7 710 11
rect 777 32 779 42
rect 784 41 786 51
rect 804 48 806 53
rect 817 48 819 53
rect 804 46 810 48
rect 804 44 806 46
rect 808 44 810 46
rect 804 42 810 44
rect 814 46 820 48
rect 814 44 816 46
rect 818 44 820 46
rect 814 42 820 44
rect 784 39 790 41
rect 784 37 786 39
rect 788 37 790 39
rect 804 38 806 42
rect 784 35 790 37
rect 784 32 786 35
rect 764 16 766 21
rect 744 7 746 11
rect 814 31 816 42
rect 824 40 826 53
rect 909 62 911 66
rect 922 64 924 69
rect 929 64 931 69
rect 953 73 978 75
rect 953 65 955 73
rect 966 65 968 69
rect 976 65 978 73
rect 986 68 988 73
rect 993 68 995 73
rect 861 53 863 56
rect 854 51 863 53
rect 871 52 873 56
rect 881 53 883 56
rect 845 43 847 51
rect 854 49 856 51
rect 858 49 863 51
rect 854 47 863 49
rect 879 51 883 53
rect 879 48 881 51
rect 861 43 863 47
rect 875 46 881 48
rect 888 47 890 56
rect 950 63 955 65
rect 950 60 952 63
rect 909 48 911 53
rect 922 48 924 53
rect 875 44 877 46
rect 879 44 881 46
rect 842 41 855 43
rect 861 41 871 43
rect 875 42 881 44
rect 842 40 844 41
rect 824 38 830 40
rect 824 36 826 38
rect 828 36 830 38
rect 824 34 830 36
rect 838 38 844 40
rect 853 38 855 41
rect 869 38 871 41
rect 879 38 881 42
rect 885 45 891 47
rect 885 43 887 45
rect 889 43 891 45
rect 885 41 891 43
rect 889 38 891 41
rect 909 46 915 48
rect 909 44 911 46
rect 913 44 915 46
rect 909 42 915 44
rect 919 46 925 48
rect 919 44 921 46
rect 923 44 925 46
rect 919 42 925 44
rect 909 38 911 42
rect 838 36 840 38
rect 842 36 844 38
rect 838 34 844 36
rect 824 31 826 34
rect 804 16 806 20
rect 814 13 816 18
rect 824 13 826 18
rect 777 7 779 11
rect 784 7 786 11
rect 869 16 871 20
rect 879 16 881 20
rect 853 7 855 11
rect 919 31 921 42
rect 929 40 931 53
rect 1024 60 1026 65
rect 966 53 968 56
rect 959 51 968 53
rect 976 52 978 56
rect 986 53 988 56
rect 950 43 952 51
rect 959 49 961 51
rect 963 49 968 51
rect 959 47 968 49
rect 984 51 988 53
rect 984 48 986 51
rect 966 43 968 47
rect 980 46 986 48
rect 993 47 995 56
rect 1034 57 1036 62
rect 1044 57 1046 62
rect 1064 62 1066 66
rect 1077 64 1079 69
rect 1084 64 1086 69
rect 1108 73 1133 75
rect 1108 65 1110 73
rect 1121 65 1123 69
rect 1131 65 1133 73
rect 1141 68 1143 73
rect 1148 68 1150 73
rect 1105 63 1110 65
rect 1105 60 1107 63
rect 1024 48 1026 51
rect 1034 48 1036 51
rect 980 44 982 46
rect 984 44 986 46
rect 947 41 960 43
rect 966 41 976 43
rect 980 42 986 44
rect 947 40 949 41
rect 929 38 935 40
rect 929 36 931 38
rect 933 36 935 38
rect 929 34 935 36
rect 943 38 949 40
rect 958 38 960 41
rect 974 38 976 41
rect 984 38 986 42
rect 990 45 996 47
rect 990 43 992 45
rect 994 43 996 45
rect 990 41 996 43
rect 994 38 996 41
rect 1024 46 1030 48
rect 1024 44 1026 46
rect 1028 44 1030 46
rect 1024 42 1030 44
rect 1034 46 1040 48
rect 1034 44 1036 46
rect 1038 44 1040 46
rect 1034 42 1040 44
rect 1024 39 1026 42
rect 943 36 945 38
rect 947 36 949 38
rect 943 34 949 36
rect 929 31 931 34
rect 909 16 911 20
rect 919 13 921 18
rect 929 13 931 18
rect 889 7 891 11
rect 974 16 976 20
rect 984 16 986 20
rect 958 7 960 11
rect 1037 32 1039 42
rect 1044 41 1046 51
rect 1064 48 1066 53
rect 1077 48 1079 53
rect 1064 46 1070 48
rect 1064 44 1066 46
rect 1068 44 1070 46
rect 1064 42 1070 44
rect 1074 46 1080 48
rect 1074 44 1076 46
rect 1078 44 1080 46
rect 1074 42 1080 44
rect 1044 39 1050 41
rect 1044 37 1046 39
rect 1048 37 1050 39
rect 1064 38 1066 42
rect 1044 35 1050 37
rect 1044 32 1046 35
rect 1024 16 1026 21
rect 994 7 996 11
rect 1074 31 1076 42
rect 1084 40 1086 53
rect 1169 62 1171 66
rect 1182 64 1184 69
rect 1189 64 1191 69
rect 1213 73 1238 75
rect 1213 65 1215 73
rect 1226 65 1228 69
rect 1236 65 1238 73
rect 1246 68 1248 73
rect 1253 68 1255 73
rect 1121 53 1123 56
rect 1114 51 1123 53
rect 1131 52 1133 56
rect 1141 53 1143 56
rect 1105 43 1107 51
rect 1114 49 1116 51
rect 1118 49 1123 51
rect 1114 47 1123 49
rect 1139 51 1143 53
rect 1139 48 1141 51
rect 1121 43 1123 47
rect 1135 46 1141 48
rect 1148 47 1150 56
rect 1210 63 1215 65
rect 1210 60 1212 63
rect 1169 48 1171 53
rect 1182 48 1184 53
rect 1135 44 1137 46
rect 1139 44 1141 46
rect 1102 41 1115 43
rect 1121 41 1131 43
rect 1135 42 1141 44
rect 1102 40 1104 41
rect 1084 38 1090 40
rect 1084 36 1086 38
rect 1088 36 1090 38
rect 1084 34 1090 36
rect 1098 38 1104 40
rect 1113 38 1115 41
rect 1129 38 1131 41
rect 1139 38 1141 42
rect 1145 45 1151 47
rect 1145 43 1147 45
rect 1149 43 1151 45
rect 1145 41 1151 43
rect 1149 38 1151 41
rect 1169 46 1175 48
rect 1169 44 1171 46
rect 1173 44 1175 46
rect 1169 42 1175 44
rect 1179 46 1185 48
rect 1179 44 1181 46
rect 1183 44 1185 46
rect 1179 42 1185 44
rect 1169 38 1171 42
rect 1098 36 1100 38
rect 1102 36 1104 38
rect 1098 34 1104 36
rect 1084 31 1086 34
rect 1064 16 1066 20
rect 1074 13 1076 18
rect 1084 13 1086 18
rect 1037 7 1039 11
rect 1044 7 1046 11
rect 1129 16 1131 20
rect 1139 16 1141 20
rect 1113 7 1115 11
rect 1179 31 1181 42
rect 1189 40 1191 53
rect 1274 60 1276 65
rect 1226 53 1228 56
rect 1219 51 1228 53
rect 1236 52 1238 56
rect 1246 53 1248 56
rect 1210 43 1212 51
rect 1219 49 1221 51
rect 1223 49 1228 51
rect 1219 47 1228 49
rect 1244 51 1248 53
rect 1244 48 1246 51
rect 1226 43 1228 47
rect 1240 46 1246 48
rect 1253 47 1255 56
rect 1284 57 1286 62
rect 1294 57 1296 62
rect 1314 62 1316 66
rect 1327 64 1329 69
rect 1334 64 1336 69
rect 1358 73 1383 75
rect 1358 65 1360 73
rect 1371 65 1373 69
rect 1381 65 1383 73
rect 1391 68 1393 73
rect 1398 68 1400 73
rect 1355 63 1360 65
rect 1355 60 1357 63
rect 1274 48 1276 51
rect 1284 48 1286 51
rect 1240 44 1242 46
rect 1244 44 1246 46
rect 1207 41 1220 43
rect 1226 41 1236 43
rect 1240 42 1246 44
rect 1207 40 1209 41
rect 1189 38 1195 40
rect 1189 36 1191 38
rect 1193 36 1195 38
rect 1189 34 1195 36
rect 1203 38 1209 40
rect 1218 38 1220 41
rect 1234 38 1236 41
rect 1244 38 1246 42
rect 1250 45 1256 47
rect 1250 43 1252 45
rect 1254 43 1256 45
rect 1250 41 1256 43
rect 1254 38 1256 41
rect 1274 46 1280 48
rect 1274 44 1276 46
rect 1278 44 1280 46
rect 1274 42 1280 44
rect 1284 46 1290 48
rect 1284 44 1286 46
rect 1288 44 1290 46
rect 1284 42 1290 44
rect 1274 39 1276 42
rect 1203 36 1205 38
rect 1207 36 1209 38
rect 1203 34 1209 36
rect 1189 31 1191 34
rect 1169 16 1171 20
rect 1179 13 1181 18
rect 1189 13 1191 18
rect 1149 7 1151 11
rect 1234 16 1236 20
rect 1244 16 1246 20
rect 1218 7 1220 11
rect 1287 32 1289 42
rect 1294 41 1296 51
rect 1314 48 1316 53
rect 1327 48 1329 53
rect 1314 46 1320 48
rect 1314 44 1316 46
rect 1318 44 1320 46
rect 1314 42 1320 44
rect 1324 46 1330 48
rect 1324 44 1326 46
rect 1328 44 1330 46
rect 1324 42 1330 44
rect 1294 39 1300 41
rect 1294 37 1296 39
rect 1298 37 1300 39
rect 1314 38 1316 42
rect 1294 35 1300 37
rect 1294 32 1296 35
rect 1274 16 1276 21
rect 1254 7 1256 11
rect 1324 31 1326 42
rect 1334 40 1336 53
rect 1419 62 1421 66
rect 1432 64 1434 69
rect 1439 64 1441 69
rect 1463 73 1488 75
rect 1463 65 1465 73
rect 1476 65 1478 69
rect 1486 65 1488 73
rect 1496 68 1498 73
rect 1503 68 1505 73
rect 1371 53 1373 56
rect 1364 51 1373 53
rect 1381 52 1383 56
rect 1391 53 1393 56
rect 1355 43 1357 51
rect 1364 49 1366 51
rect 1368 49 1373 51
rect 1364 47 1373 49
rect 1389 51 1393 53
rect 1389 48 1391 51
rect 1371 43 1373 47
rect 1385 46 1391 48
rect 1398 47 1400 56
rect 1460 63 1465 65
rect 1460 60 1462 63
rect 1419 48 1421 53
rect 1432 48 1434 53
rect 1385 44 1387 46
rect 1389 44 1391 46
rect 1352 41 1365 43
rect 1371 41 1381 43
rect 1385 42 1391 44
rect 1352 40 1354 41
rect 1334 38 1340 40
rect 1334 36 1336 38
rect 1338 36 1340 38
rect 1334 34 1340 36
rect 1348 38 1354 40
rect 1363 38 1365 41
rect 1379 38 1381 41
rect 1389 38 1391 42
rect 1395 45 1401 47
rect 1395 43 1397 45
rect 1399 43 1401 45
rect 1395 41 1401 43
rect 1399 38 1401 41
rect 1419 46 1425 48
rect 1419 44 1421 46
rect 1423 44 1425 46
rect 1419 42 1425 44
rect 1429 46 1435 48
rect 1429 44 1431 46
rect 1433 44 1435 46
rect 1429 42 1435 44
rect 1419 38 1421 42
rect 1348 36 1350 38
rect 1352 36 1354 38
rect 1348 34 1354 36
rect 1334 31 1336 34
rect 1314 16 1316 20
rect 1324 13 1326 18
rect 1334 13 1336 18
rect 1287 7 1289 11
rect 1294 7 1296 11
rect 1379 16 1381 20
rect 1389 16 1391 20
rect 1363 7 1365 11
rect 1429 31 1431 42
rect 1439 40 1441 53
rect 1524 60 1526 65
rect 1476 53 1478 56
rect 1469 51 1478 53
rect 1486 52 1488 56
rect 1496 53 1498 56
rect 1460 43 1462 51
rect 1469 49 1471 51
rect 1473 49 1478 51
rect 1469 47 1478 49
rect 1494 51 1498 53
rect 1494 48 1496 51
rect 1476 43 1478 47
rect 1490 46 1496 48
rect 1503 47 1505 56
rect 1534 57 1536 62
rect 1544 57 1546 62
rect 1564 62 1566 66
rect 1577 64 1579 69
rect 1584 64 1586 69
rect 1608 73 1633 75
rect 1608 65 1610 73
rect 1621 65 1623 69
rect 1631 65 1633 73
rect 1641 68 1643 73
rect 1648 68 1650 73
rect 1605 63 1610 65
rect 1605 60 1607 63
rect 1524 48 1526 51
rect 1534 48 1536 51
rect 1490 44 1492 46
rect 1494 44 1496 46
rect 1457 41 1470 43
rect 1476 41 1486 43
rect 1490 42 1496 44
rect 1457 40 1459 41
rect 1439 38 1445 40
rect 1439 36 1441 38
rect 1443 36 1445 38
rect 1439 34 1445 36
rect 1453 38 1459 40
rect 1468 38 1470 41
rect 1484 38 1486 41
rect 1494 38 1496 42
rect 1500 45 1506 47
rect 1500 43 1502 45
rect 1504 43 1506 45
rect 1500 41 1506 43
rect 1504 38 1506 41
rect 1524 46 1530 48
rect 1524 44 1526 46
rect 1528 44 1530 46
rect 1524 42 1530 44
rect 1534 46 1540 48
rect 1534 44 1536 46
rect 1538 44 1540 46
rect 1534 42 1540 44
rect 1524 39 1526 42
rect 1453 36 1455 38
rect 1457 36 1459 38
rect 1453 34 1459 36
rect 1439 31 1441 34
rect 1419 16 1421 20
rect 1429 13 1431 18
rect 1439 13 1441 18
rect 1399 7 1401 11
rect 1484 16 1486 20
rect 1494 16 1496 20
rect 1468 7 1470 11
rect 1537 32 1539 42
rect 1544 41 1546 51
rect 1564 48 1566 53
rect 1577 48 1579 53
rect 1564 46 1570 48
rect 1564 44 1566 46
rect 1568 44 1570 46
rect 1564 42 1570 44
rect 1574 46 1580 48
rect 1574 44 1576 46
rect 1578 44 1580 46
rect 1574 42 1580 44
rect 1544 39 1550 41
rect 1544 37 1546 39
rect 1548 37 1550 39
rect 1564 38 1566 42
rect 1544 35 1550 37
rect 1544 32 1546 35
rect 1524 16 1526 21
rect 1504 7 1506 11
rect 1574 31 1576 42
rect 1584 40 1586 53
rect 1669 62 1671 66
rect 1682 64 1684 69
rect 1689 64 1691 69
rect 1713 73 1738 75
rect 1713 65 1715 73
rect 1726 65 1728 69
rect 1736 65 1738 73
rect 1746 68 1748 73
rect 1753 68 1755 73
rect 1621 53 1623 56
rect 1614 51 1623 53
rect 1631 52 1633 56
rect 1641 53 1643 56
rect 1605 43 1607 51
rect 1614 49 1616 51
rect 1618 49 1623 51
rect 1614 47 1623 49
rect 1639 51 1643 53
rect 1639 48 1641 51
rect 1621 43 1623 47
rect 1635 46 1641 48
rect 1648 47 1650 56
rect 1710 63 1715 65
rect 1710 60 1712 63
rect 1669 48 1671 53
rect 1682 48 1684 53
rect 1635 44 1637 46
rect 1639 44 1641 46
rect 1602 41 1615 43
rect 1621 41 1631 43
rect 1635 42 1641 44
rect 1602 40 1604 41
rect 1584 38 1590 40
rect 1584 36 1586 38
rect 1588 36 1590 38
rect 1584 34 1590 36
rect 1598 38 1604 40
rect 1613 38 1615 41
rect 1629 38 1631 41
rect 1639 38 1641 42
rect 1645 45 1651 47
rect 1645 43 1647 45
rect 1649 43 1651 45
rect 1645 41 1651 43
rect 1649 38 1651 41
rect 1669 46 1675 48
rect 1669 44 1671 46
rect 1673 44 1675 46
rect 1669 42 1675 44
rect 1679 46 1685 48
rect 1679 44 1681 46
rect 1683 44 1685 46
rect 1679 42 1685 44
rect 1669 38 1671 42
rect 1598 36 1600 38
rect 1602 36 1604 38
rect 1598 34 1604 36
rect 1584 31 1586 34
rect 1564 16 1566 20
rect 1574 13 1576 18
rect 1584 13 1586 18
rect 1537 7 1539 11
rect 1544 7 1546 11
rect 1629 16 1631 20
rect 1639 16 1641 20
rect 1613 7 1615 11
rect 1679 31 1681 42
rect 1689 40 1691 53
rect 1774 60 1776 65
rect 1726 53 1728 56
rect 1719 51 1728 53
rect 1736 52 1738 56
rect 1746 53 1748 56
rect 1710 43 1712 51
rect 1719 49 1721 51
rect 1723 49 1728 51
rect 1719 47 1728 49
rect 1744 51 1748 53
rect 1744 48 1746 51
rect 1726 43 1728 47
rect 1740 46 1746 48
rect 1753 47 1755 56
rect 1784 57 1786 62
rect 1794 57 1796 62
rect 1814 62 1816 66
rect 1827 64 1829 69
rect 1834 64 1836 69
rect 1858 73 1883 75
rect 1858 65 1860 73
rect 1871 65 1873 69
rect 1881 65 1883 73
rect 1891 68 1893 73
rect 1898 68 1900 73
rect 1855 63 1860 65
rect 1855 60 1857 63
rect 1774 48 1776 51
rect 1784 48 1786 51
rect 1740 44 1742 46
rect 1744 44 1746 46
rect 1707 41 1720 43
rect 1726 41 1736 43
rect 1740 42 1746 44
rect 1707 40 1709 41
rect 1689 38 1695 40
rect 1689 36 1691 38
rect 1693 36 1695 38
rect 1689 34 1695 36
rect 1703 38 1709 40
rect 1718 38 1720 41
rect 1734 38 1736 41
rect 1744 38 1746 42
rect 1750 45 1756 47
rect 1750 43 1752 45
rect 1754 43 1756 45
rect 1750 41 1756 43
rect 1754 38 1756 41
rect 1774 46 1780 48
rect 1774 44 1776 46
rect 1778 44 1780 46
rect 1774 42 1780 44
rect 1784 46 1790 48
rect 1784 44 1786 46
rect 1788 44 1790 46
rect 1784 42 1790 44
rect 1774 39 1776 42
rect 1703 36 1705 38
rect 1707 36 1709 38
rect 1703 34 1709 36
rect 1689 31 1691 34
rect 1669 16 1671 20
rect 1679 13 1681 18
rect 1689 13 1691 18
rect 1649 7 1651 11
rect 1734 16 1736 20
rect 1744 16 1746 20
rect 1718 7 1720 11
rect 1787 32 1789 42
rect 1794 41 1796 51
rect 1814 48 1816 53
rect 1827 48 1829 53
rect 1814 46 1820 48
rect 1814 44 1816 46
rect 1818 44 1820 46
rect 1814 42 1820 44
rect 1824 46 1830 48
rect 1824 44 1826 46
rect 1828 44 1830 46
rect 1824 42 1830 44
rect 1794 39 1800 41
rect 1794 37 1796 39
rect 1798 37 1800 39
rect 1814 38 1816 42
rect 1794 35 1800 37
rect 1794 32 1796 35
rect 1774 16 1776 21
rect 1754 7 1756 11
rect 1824 31 1826 42
rect 1834 40 1836 53
rect 1919 62 1921 66
rect 1932 64 1934 69
rect 1939 64 1941 69
rect 1963 73 1988 75
rect 1963 65 1965 73
rect 1976 65 1978 69
rect 1986 65 1988 73
rect 1996 68 1998 73
rect 2003 68 2005 73
rect 1871 53 1873 56
rect 1864 51 1873 53
rect 1881 52 1883 56
rect 1891 53 1893 56
rect 1855 43 1857 51
rect 1864 49 1866 51
rect 1868 49 1873 51
rect 1864 47 1873 49
rect 1889 51 1893 53
rect 1889 48 1891 51
rect 1871 43 1873 47
rect 1885 46 1891 48
rect 1898 47 1900 56
rect 1960 63 1965 65
rect 1960 60 1962 63
rect 1919 48 1921 53
rect 1932 48 1934 53
rect 1885 44 1887 46
rect 1889 44 1891 46
rect 1852 41 1865 43
rect 1871 41 1881 43
rect 1885 42 1891 44
rect 1852 40 1854 41
rect 1834 38 1840 40
rect 1834 36 1836 38
rect 1838 36 1840 38
rect 1834 34 1840 36
rect 1848 38 1854 40
rect 1863 38 1865 41
rect 1879 38 1881 41
rect 1889 38 1891 42
rect 1895 45 1901 47
rect 1895 43 1897 45
rect 1899 43 1901 45
rect 1895 41 1901 43
rect 1899 38 1901 41
rect 1919 46 1925 48
rect 1919 44 1921 46
rect 1923 44 1925 46
rect 1919 42 1925 44
rect 1929 46 1935 48
rect 1929 44 1931 46
rect 1933 44 1935 46
rect 1929 42 1935 44
rect 1919 38 1921 42
rect 1848 36 1850 38
rect 1852 36 1854 38
rect 1848 34 1854 36
rect 1834 31 1836 34
rect 1814 16 1816 20
rect 1824 13 1826 18
rect 1834 13 1836 18
rect 1787 7 1789 11
rect 1794 7 1796 11
rect 1879 16 1881 20
rect 1889 16 1891 20
rect 1863 7 1865 11
rect 1929 31 1931 42
rect 1939 40 1941 53
rect 1976 53 1978 56
rect 1969 51 1978 53
rect 1986 52 1988 56
rect 1996 53 1998 56
rect 1960 43 1962 51
rect 1969 49 1971 51
rect 1973 49 1978 51
rect 1969 47 1978 49
rect 1994 51 1998 53
rect 1994 48 1996 51
rect 1976 43 1978 47
rect 1990 46 1996 48
rect 2003 47 2005 56
rect 1990 44 1992 46
rect 1994 44 1996 46
rect 1957 41 1970 43
rect 1976 41 1986 43
rect 1990 42 1996 44
rect 1957 40 1959 41
rect 1939 38 1945 40
rect 1939 36 1941 38
rect 1943 36 1945 38
rect 1939 34 1945 36
rect 1953 38 1959 40
rect 1968 38 1970 41
rect 1984 38 1986 41
rect 1994 38 1996 42
rect 2000 45 2006 47
rect 2000 43 2002 45
rect 2004 43 2006 45
rect 2000 41 2006 43
rect 2004 38 2006 41
rect 1953 36 1955 38
rect 1957 36 1959 38
rect 1953 34 1959 36
rect 1939 31 1941 34
rect 1919 16 1921 20
rect 1929 13 1931 18
rect 1939 13 1941 18
rect 1899 7 1901 11
rect 1984 16 1986 20
rect 1994 16 1996 20
rect 1968 7 1970 11
rect 2004 7 2006 11
<< ndif >>
rect 51 226 58 228
rect 51 224 54 226
rect 56 224 58 226
rect 51 218 58 224
rect 91 226 98 228
rect 91 224 94 226
rect 96 224 98 226
rect 33 216 40 218
rect 33 214 35 216
rect 37 214 40 216
rect 33 212 40 214
rect 35 207 40 212
rect 42 207 47 218
rect 49 216 58 218
rect 91 218 98 224
rect 120 226 126 228
rect 120 224 122 226
rect 124 224 126 226
rect 120 222 126 224
rect 73 216 80 218
rect 49 207 60 216
rect 62 214 69 216
rect 62 212 65 214
rect 67 212 69 214
rect 73 214 75 216
rect 77 214 80 216
rect 73 212 80 214
rect 62 210 69 212
rect 62 207 67 210
rect 75 207 80 212
rect 82 207 87 218
rect 89 216 98 218
rect 89 207 100 216
rect 102 214 109 216
rect 102 212 105 214
rect 107 212 109 214
rect 102 210 109 212
rect 120 210 128 222
rect 130 210 135 222
rect 137 219 142 222
rect 203 226 210 228
rect 203 224 206 226
rect 208 224 210 226
rect 137 216 145 219
rect 137 214 140 216
rect 142 214 145 216
rect 137 210 145 214
rect 147 214 155 219
rect 147 212 150 214
rect 152 212 155 214
rect 147 210 155 212
rect 157 217 166 219
rect 203 218 210 224
rect 374 225 381 227
rect 374 223 376 225
rect 378 223 381 225
rect 157 215 162 217
rect 164 215 166 217
rect 157 214 166 215
rect 185 216 192 218
rect 185 214 187 216
rect 189 214 192 216
rect 157 210 171 214
rect 102 207 107 210
rect 166 205 171 210
rect 173 211 178 214
rect 185 212 192 214
rect 173 209 180 211
rect 173 207 176 209
rect 178 207 180 209
rect 187 207 192 212
rect 194 207 199 218
rect 201 216 210 218
rect 201 207 212 216
rect 214 214 221 216
rect 374 217 381 223
rect 421 225 428 227
rect 421 223 424 225
rect 426 223 428 225
rect 421 217 428 223
rect 454 225 461 227
rect 454 223 456 225
rect 458 223 461 225
rect 374 215 383 217
rect 214 212 217 214
rect 219 212 221 214
rect 214 210 221 212
rect 363 213 370 215
rect 363 211 365 213
rect 367 211 370 213
rect 214 207 219 210
rect 363 209 370 211
rect 173 205 180 207
rect 365 206 370 209
rect 372 206 383 215
rect 385 206 390 217
rect 392 215 399 217
rect 392 213 395 215
rect 397 213 399 215
rect 392 211 399 213
rect 403 215 410 217
rect 403 213 405 215
rect 407 213 410 215
rect 403 211 410 213
rect 392 206 397 211
rect 405 206 410 211
rect 412 206 417 217
rect 419 215 428 217
rect 454 217 461 223
rect 538 225 544 227
rect 538 223 540 225
rect 542 223 544 225
rect 538 221 544 223
rect 579 225 586 227
rect 579 223 581 225
rect 583 223 586 225
rect 522 218 527 221
rect 454 215 463 217
rect 419 206 430 215
rect 432 213 439 215
rect 432 211 435 213
rect 437 211 439 213
rect 432 209 439 211
rect 443 213 450 215
rect 443 211 445 213
rect 447 211 450 213
rect 443 209 450 211
rect 432 206 437 209
rect 445 206 450 209
rect 452 206 463 215
rect 465 206 470 217
rect 472 215 479 217
rect 472 213 475 215
rect 477 213 479 215
rect 498 216 507 218
rect 498 214 500 216
rect 502 214 507 216
rect 498 213 507 214
rect 472 211 479 213
rect 472 206 477 211
rect 486 210 491 213
rect 484 208 491 210
rect 484 206 486 208
rect 488 206 491 208
rect 484 204 491 206
rect 493 209 507 213
rect 509 213 517 218
rect 509 211 512 213
rect 514 211 517 213
rect 509 209 517 211
rect 519 215 527 218
rect 519 213 522 215
rect 524 213 527 215
rect 519 209 527 213
rect 529 209 534 221
rect 536 209 544 221
rect 579 217 586 223
rect 626 225 633 227
rect 626 223 629 225
rect 631 223 633 225
rect 626 217 633 223
rect 659 225 666 227
rect 659 223 661 225
rect 663 223 666 225
rect 579 215 588 217
rect 568 213 575 215
rect 568 211 570 213
rect 572 211 575 213
rect 568 209 575 211
rect 493 204 498 209
rect 570 206 575 209
rect 577 206 588 215
rect 590 206 595 217
rect 597 215 604 217
rect 597 213 600 215
rect 602 213 604 215
rect 597 211 604 213
rect 608 215 615 217
rect 608 213 610 215
rect 612 213 615 215
rect 608 211 615 213
rect 597 206 602 211
rect 610 206 615 211
rect 617 206 622 217
rect 624 215 633 217
rect 659 217 666 223
rect 743 225 749 227
rect 743 223 745 225
rect 747 223 749 225
rect 1841 226 1848 228
rect 1841 224 1844 226
rect 1846 224 1848 226
rect 743 221 749 223
rect 727 218 732 221
rect 659 215 668 217
rect 624 206 635 215
rect 637 213 644 215
rect 637 211 640 213
rect 642 211 644 213
rect 637 209 644 211
rect 648 213 655 215
rect 648 211 650 213
rect 652 211 655 213
rect 648 209 655 211
rect 637 206 642 209
rect 650 206 655 209
rect 657 206 668 215
rect 670 206 675 217
rect 677 215 684 217
rect 677 213 680 215
rect 682 213 684 215
rect 703 216 712 218
rect 703 214 705 216
rect 707 214 712 216
rect 703 213 712 214
rect 677 211 684 213
rect 677 206 682 211
rect 691 210 696 213
rect 689 208 696 210
rect 689 206 691 208
rect 693 206 696 208
rect 689 204 696 206
rect 698 209 712 213
rect 714 213 722 218
rect 714 211 717 213
rect 719 211 722 213
rect 714 209 722 211
rect 724 215 732 218
rect 724 213 727 215
rect 729 213 732 215
rect 724 209 732 213
rect 734 209 739 221
rect 741 209 749 221
rect 1841 218 1848 224
rect 1881 226 1888 228
rect 1881 224 1884 226
rect 1886 224 1888 226
rect 1823 216 1830 218
rect 1823 214 1825 216
rect 1827 214 1830 216
rect 1823 212 1830 214
rect 698 204 703 209
rect 1825 207 1830 212
rect 1832 207 1837 218
rect 1839 216 1848 218
rect 1881 218 1888 224
rect 1910 226 1916 228
rect 1910 224 1912 226
rect 1914 224 1916 226
rect 1910 222 1916 224
rect 1863 216 1870 218
rect 1839 207 1850 216
rect 1852 214 1859 216
rect 1852 212 1855 214
rect 1857 212 1859 214
rect 1863 214 1865 216
rect 1867 214 1870 216
rect 1863 212 1870 214
rect 1852 210 1859 212
rect 1852 207 1857 210
rect 1865 207 1870 212
rect 1872 207 1877 218
rect 1879 216 1888 218
rect 1879 207 1890 216
rect 1892 214 1899 216
rect 1892 212 1895 214
rect 1897 212 1899 214
rect 1892 210 1899 212
rect 1910 210 1918 222
rect 1920 210 1925 222
rect 1927 219 1932 222
rect 1993 226 2000 228
rect 1993 224 1996 226
rect 1998 224 2000 226
rect 1927 216 1935 219
rect 1927 214 1930 216
rect 1932 214 1935 216
rect 1927 210 1935 214
rect 1937 214 1945 219
rect 1937 212 1940 214
rect 1942 212 1945 214
rect 1937 210 1945 212
rect 1947 217 1956 219
rect 1993 218 2000 224
rect 1947 215 1952 217
rect 1954 215 1956 217
rect 1947 214 1956 215
rect 1975 216 1982 218
rect 1975 214 1977 216
rect 1979 214 1982 216
rect 1947 210 1961 214
rect 1892 207 1897 210
rect 1956 205 1961 210
rect 1963 211 1968 214
rect 1975 212 1982 214
rect 1963 209 1970 211
rect 1963 207 1966 209
rect 1968 207 1970 209
rect 1977 207 1982 212
rect 1984 207 1989 218
rect 1991 216 2000 218
rect 1991 207 2002 216
rect 2004 214 2011 216
rect 2004 212 2007 214
rect 2009 212 2011 214
rect 2004 210 2011 212
rect 2004 207 2009 210
rect 1963 205 1970 207
rect 154 111 161 113
rect 35 108 40 111
rect 33 106 40 108
rect 33 104 35 106
rect 37 104 40 106
rect 33 102 40 104
rect 42 102 53 111
rect 44 100 53 102
rect 55 100 60 111
rect 62 106 67 111
rect 75 106 80 111
rect 62 104 69 106
rect 62 102 65 104
rect 67 102 69 104
rect 62 100 69 102
rect 73 104 80 106
rect 73 102 75 104
rect 77 102 80 104
rect 73 100 80 102
rect 82 100 87 111
rect 89 102 100 111
rect 102 108 107 111
rect 115 108 120 111
rect 102 106 109 108
rect 102 104 105 106
rect 107 104 109 106
rect 102 102 109 104
rect 113 106 120 108
rect 113 104 115 106
rect 117 104 120 106
rect 113 102 120 104
rect 122 102 133 111
rect 89 100 98 102
rect 44 94 51 100
rect 44 92 46 94
rect 48 92 51 94
rect 44 90 51 92
rect 91 94 98 100
rect 124 100 133 102
rect 135 100 140 111
rect 142 106 147 111
rect 154 109 156 111
rect 158 109 161 111
rect 154 107 161 109
rect 142 104 149 106
rect 156 104 161 107
rect 163 108 168 113
rect 278 111 285 113
rect 239 108 244 111
rect 163 104 177 108
rect 142 102 145 104
rect 147 102 149 104
rect 142 100 149 102
rect 168 103 177 104
rect 168 101 170 103
rect 172 101 177 103
rect 91 92 94 94
rect 96 92 98 94
rect 91 90 98 92
rect 124 94 131 100
rect 168 99 177 101
rect 179 106 187 108
rect 179 104 182 106
rect 184 104 187 106
rect 179 99 187 104
rect 189 104 197 108
rect 189 102 192 104
rect 194 102 197 104
rect 189 99 197 102
rect 124 92 126 94
rect 128 92 131 94
rect 124 90 131 92
rect 192 96 197 99
rect 199 96 204 108
rect 206 96 214 108
rect 237 106 244 108
rect 237 104 239 106
rect 241 104 244 106
rect 237 102 244 104
rect 246 102 257 111
rect 248 100 257 102
rect 259 100 264 111
rect 266 106 271 111
rect 278 109 280 111
rect 282 109 285 111
rect 278 107 285 109
rect 266 104 273 106
rect 280 104 285 107
rect 287 108 292 113
rect 287 104 301 108
rect 266 102 269 104
rect 271 102 273 104
rect 266 100 273 102
rect 292 103 301 104
rect 292 101 294 103
rect 296 101 301 103
rect 208 94 214 96
rect 208 92 210 94
rect 212 92 214 94
rect 208 90 214 92
rect 248 94 255 100
rect 292 99 301 101
rect 303 106 311 108
rect 303 104 306 106
rect 308 104 311 106
rect 303 99 311 104
rect 313 104 321 108
rect 313 102 316 104
rect 318 102 321 104
rect 313 99 321 102
rect 248 92 250 94
rect 252 92 255 94
rect 248 90 255 92
rect 316 96 321 99
rect 323 96 328 108
rect 330 96 338 108
rect 365 105 370 110
rect 363 103 370 105
rect 363 101 365 103
rect 367 101 370 103
rect 363 99 370 101
rect 372 99 377 110
rect 379 101 390 110
rect 392 107 397 110
rect 392 105 399 107
rect 405 105 410 110
rect 392 103 395 105
rect 397 103 399 105
rect 392 101 399 103
rect 403 103 410 105
rect 403 101 405 103
rect 407 101 410 103
rect 379 99 388 101
rect 332 94 338 96
rect 332 92 334 94
rect 336 92 338 94
rect 332 90 338 92
rect 381 93 388 99
rect 403 99 410 101
rect 412 99 417 110
rect 419 101 430 110
rect 432 107 437 110
rect 496 107 501 112
rect 432 105 439 107
rect 432 103 435 105
rect 437 103 439 105
rect 432 101 439 103
rect 419 99 428 101
rect 381 91 384 93
rect 386 91 388 93
rect 381 89 388 91
rect 421 93 428 99
rect 450 95 458 107
rect 460 95 465 107
rect 467 103 475 107
rect 467 101 470 103
rect 472 101 475 103
rect 467 98 475 101
rect 477 105 485 107
rect 477 103 480 105
rect 482 103 485 105
rect 477 98 485 103
rect 487 103 501 107
rect 503 110 510 112
rect 503 108 506 110
rect 508 108 510 110
rect 503 106 510 108
rect 503 103 508 106
rect 517 105 522 110
rect 515 103 522 105
rect 487 102 496 103
rect 487 100 492 102
rect 494 100 496 102
rect 487 98 496 100
rect 515 101 517 103
rect 519 101 522 103
rect 515 99 522 101
rect 524 99 529 110
rect 531 101 542 110
rect 544 107 549 110
rect 544 105 551 107
rect 570 105 575 110
rect 544 103 547 105
rect 549 103 551 105
rect 544 101 551 103
rect 568 103 575 105
rect 568 101 570 103
rect 572 101 575 103
rect 531 99 540 101
rect 467 95 472 98
rect 421 91 424 93
rect 426 91 428 93
rect 421 89 428 91
rect 450 93 456 95
rect 450 91 452 93
rect 454 91 456 93
rect 450 89 456 91
rect 533 93 540 99
rect 568 99 575 101
rect 577 99 582 110
rect 584 101 595 110
rect 597 107 602 110
rect 597 105 604 107
rect 610 105 615 110
rect 597 103 600 105
rect 602 103 604 105
rect 597 101 604 103
rect 608 103 615 105
rect 608 101 610 103
rect 612 101 615 103
rect 584 99 593 101
rect 533 91 536 93
rect 538 91 540 93
rect 533 89 540 91
rect 586 93 593 99
rect 608 99 615 101
rect 617 99 622 110
rect 624 101 635 110
rect 637 107 642 110
rect 701 107 706 112
rect 637 105 644 107
rect 637 103 640 105
rect 642 103 644 105
rect 637 101 644 103
rect 624 99 633 101
rect 586 91 589 93
rect 591 91 593 93
rect 586 89 593 91
rect 626 93 633 99
rect 655 95 663 107
rect 665 95 670 107
rect 672 103 680 107
rect 672 101 675 103
rect 677 101 680 103
rect 672 98 680 101
rect 682 105 690 107
rect 682 103 685 105
rect 687 103 690 105
rect 682 98 690 103
rect 692 103 706 107
rect 708 110 715 112
rect 775 111 782 113
rect 708 108 711 110
rect 713 108 715 110
rect 708 106 715 108
rect 708 103 713 106
rect 722 105 727 110
rect 720 103 727 105
rect 692 102 701 103
rect 692 100 697 102
rect 699 100 701 102
rect 692 98 701 100
rect 720 101 722 103
rect 724 101 727 103
rect 720 99 727 101
rect 729 99 734 110
rect 736 101 747 110
rect 749 107 754 110
rect 775 109 777 111
rect 779 109 782 111
rect 775 107 782 109
rect 749 105 756 107
rect 749 103 752 105
rect 754 103 756 105
rect 777 104 782 107
rect 784 107 792 113
rect 794 111 802 113
rect 794 109 797 111
rect 799 109 802 111
rect 794 107 802 109
rect 804 107 811 113
rect 856 111 863 113
rect 817 108 822 111
rect 784 104 790 107
rect 749 101 756 103
rect 736 99 745 101
rect 672 95 677 98
rect 626 91 629 93
rect 631 91 633 93
rect 626 89 633 91
rect 655 93 661 95
rect 655 91 657 93
rect 659 91 661 93
rect 655 89 661 91
rect 738 93 745 99
rect 786 100 790 104
rect 806 100 811 107
rect 815 106 822 108
rect 815 104 817 106
rect 819 104 822 106
rect 815 102 822 104
rect 824 102 835 111
rect 786 98 792 100
rect 786 96 788 98
rect 790 96 792 98
rect 738 91 741 93
rect 743 91 745 93
rect 738 89 745 91
rect 786 94 792 96
rect 805 98 811 100
rect 826 100 835 102
rect 837 100 842 111
rect 844 106 849 111
rect 856 109 858 111
rect 860 109 863 111
rect 856 107 863 109
rect 844 104 851 106
rect 858 104 863 107
rect 865 108 870 113
rect 961 111 968 113
rect 922 108 927 111
rect 865 104 879 108
rect 844 102 847 104
rect 849 102 851 104
rect 844 100 851 102
rect 870 103 879 104
rect 870 101 872 103
rect 874 101 879 103
rect 805 96 807 98
rect 809 96 811 98
rect 805 94 811 96
rect 826 94 833 100
rect 870 99 879 101
rect 881 106 889 108
rect 881 104 884 106
rect 886 104 889 106
rect 881 99 889 104
rect 891 104 899 108
rect 891 102 894 104
rect 896 102 899 104
rect 891 99 899 102
rect 826 92 828 94
rect 830 92 833 94
rect 826 90 833 92
rect 894 96 899 99
rect 901 96 906 108
rect 908 96 916 108
rect 920 106 927 108
rect 920 104 922 106
rect 924 104 927 106
rect 920 102 927 104
rect 929 102 940 111
rect 931 100 940 102
rect 942 100 947 111
rect 949 106 954 111
rect 961 109 963 111
rect 965 109 968 111
rect 961 107 968 109
rect 949 104 956 106
rect 963 104 968 107
rect 970 108 975 113
rect 1025 111 1032 113
rect 1025 109 1027 111
rect 1029 109 1032 111
rect 970 104 984 108
rect 949 102 952 104
rect 954 102 956 104
rect 949 100 956 102
rect 975 103 984 104
rect 975 101 977 103
rect 979 101 984 103
rect 910 94 916 96
rect 910 92 912 94
rect 914 92 916 94
rect 910 90 916 92
rect 931 94 938 100
rect 975 99 984 101
rect 986 106 994 108
rect 986 104 989 106
rect 991 104 994 106
rect 986 99 994 104
rect 996 104 1004 108
rect 996 102 999 104
rect 1001 102 1004 104
rect 996 99 1004 102
rect 931 92 933 94
rect 935 92 938 94
rect 931 90 938 92
rect 999 96 1004 99
rect 1006 96 1011 108
rect 1013 96 1021 108
rect 1025 107 1032 109
rect 1027 104 1032 107
rect 1034 107 1042 113
rect 1044 111 1052 113
rect 1044 109 1047 111
rect 1049 109 1052 111
rect 1044 107 1052 109
rect 1054 107 1061 113
rect 1106 111 1113 113
rect 1067 108 1072 111
rect 1034 104 1040 107
rect 1036 100 1040 104
rect 1056 100 1061 107
rect 1065 106 1072 108
rect 1065 104 1067 106
rect 1069 104 1072 106
rect 1065 102 1072 104
rect 1074 102 1085 111
rect 1036 98 1042 100
rect 1036 96 1038 98
rect 1040 96 1042 98
rect 1015 94 1021 96
rect 1015 92 1017 94
rect 1019 92 1021 94
rect 1015 90 1021 92
rect 1036 94 1042 96
rect 1055 98 1061 100
rect 1076 100 1085 102
rect 1087 100 1092 111
rect 1094 106 1099 111
rect 1106 109 1108 111
rect 1110 109 1113 111
rect 1106 107 1113 109
rect 1094 104 1101 106
rect 1108 104 1113 107
rect 1115 108 1120 113
rect 1211 111 1218 113
rect 1172 108 1177 111
rect 1115 104 1129 108
rect 1094 102 1097 104
rect 1099 102 1101 104
rect 1094 100 1101 102
rect 1120 103 1129 104
rect 1120 101 1122 103
rect 1124 101 1129 103
rect 1055 96 1057 98
rect 1059 96 1061 98
rect 1055 94 1061 96
rect 1076 94 1083 100
rect 1120 99 1129 101
rect 1131 106 1139 108
rect 1131 104 1134 106
rect 1136 104 1139 106
rect 1131 99 1139 104
rect 1141 104 1149 108
rect 1141 102 1144 104
rect 1146 102 1149 104
rect 1141 99 1149 102
rect 1076 92 1078 94
rect 1080 92 1083 94
rect 1076 90 1083 92
rect 1144 96 1149 99
rect 1151 96 1156 108
rect 1158 96 1166 108
rect 1170 106 1177 108
rect 1170 104 1172 106
rect 1174 104 1177 106
rect 1170 102 1177 104
rect 1179 102 1190 111
rect 1181 100 1190 102
rect 1192 100 1197 111
rect 1199 106 1204 111
rect 1211 109 1213 111
rect 1215 109 1218 111
rect 1211 107 1218 109
rect 1199 104 1206 106
rect 1213 104 1218 107
rect 1220 108 1225 113
rect 1275 111 1282 113
rect 1275 109 1277 111
rect 1279 109 1282 111
rect 1220 104 1234 108
rect 1199 102 1202 104
rect 1204 102 1206 104
rect 1199 100 1206 102
rect 1225 103 1234 104
rect 1225 101 1227 103
rect 1229 101 1234 103
rect 1160 94 1166 96
rect 1160 92 1162 94
rect 1164 92 1166 94
rect 1160 90 1166 92
rect 1181 94 1188 100
rect 1225 99 1234 101
rect 1236 106 1244 108
rect 1236 104 1239 106
rect 1241 104 1244 106
rect 1236 99 1244 104
rect 1246 104 1254 108
rect 1246 102 1249 104
rect 1251 102 1254 104
rect 1246 99 1254 102
rect 1181 92 1183 94
rect 1185 92 1188 94
rect 1181 90 1188 92
rect 1249 96 1254 99
rect 1256 96 1261 108
rect 1263 96 1271 108
rect 1275 107 1282 109
rect 1277 104 1282 107
rect 1284 107 1292 113
rect 1294 111 1302 113
rect 1294 109 1297 111
rect 1299 109 1302 111
rect 1294 107 1302 109
rect 1304 107 1311 113
rect 1356 111 1363 113
rect 1317 108 1322 111
rect 1284 104 1290 107
rect 1286 100 1290 104
rect 1306 100 1311 107
rect 1315 106 1322 108
rect 1315 104 1317 106
rect 1319 104 1322 106
rect 1315 102 1322 104
rect 1324 102 1335 111
rect 1286 98 1292 100
rect 1286 96 1288 98
rect 1290 96 1292 98
rect 1265 94 1271 96
rect 1265 92 1267 94
rect 1269 92 1271 94
rect 1265 90 1271 92
rect 1286 94 1292 96
rect 1305 98 1311 100
rect 1326 100 1335 102
rect 1337 100 1342 111
rect 1344 106 1349 111
rect 1356 109 1358 111
rect 1360 109 1363 111
rect 1356 107 1363 109
rect 1344 104 1351 106
rect 1358 104 1363 107
rect 1365 108 1370 113
rect 1461 111 1468 113
rect 1422 108 1427 111
rect 1365 104 1379 108
rect 1344 102 1347 104
rect 1349 102 1351 104
rect 1344 100 1351 102
rect 1370 103 1379 104
rect 1370 101 1372 103
rect 1374 101 1379 103
rect 1305 96 1307 98
rect 1309 96 1311 98
rect 1305 94 1311 96
rect 1326 94 1333 100
rect 1370 99 1379 101
rect 1381 106 1389 108
rect 1381 104 1384 106
rect 1386 104 1389 106
rect 1381 99 1389 104
rect 1391 104 1399 108
rect 1391 102 1394 104
rect 1396 102 1399 104
rect 1391 99 1399 102
rect 1326 92 1328 94
rect 1330 92 1333 94
rect 1326 90 1333 92
rect 1394 96 1399 99
rect 1401 96 1406 108
rect 1408 96 1416 108
rect 1420 106 1427 108
rect 1420 104 1422 106
rect 1424 104 1427 106
rect 1420 102 1427 104
rect 1429 102 1440 111
rect 1431 100 1440 102
rect 1442 100 1447 111
rect 1449 106 1454 111
rect 1461 109 1463 111
rect 1465 109 1468 111
rect 1461 107 1468 109
rect 1449 104 1456 106
rect 1463 104 1468 107
rect 1470 108 1475 113
rect 1525 111 1532 113
rect 1525 109 1527 111
rect 1529 109 1532 111
rect 1470 104 1484 108
rect 1449 102 1452 104
rect 1454 102 1456 104
rect 1449 100 1456 102
rect 1475 103 1484 104
rect 1475 101 1477 103
rect 1479 101 1484 103
rect 1410 94 1416 96
rect 1410 92 1412 94
rect 1414 92 1416 94
rect 1410 90 1416 92
rect 1431 94 1438 100
rect 1475 99 1484 101
rect 1486 106 1494 108
rect 1486 104 1489 106
rect 1491 104 1494 106
rect 1486 99 1494 104
rect 1496 104 1504 108
rect 1496 102 1499 104
rect 1501 102 1504 104
rect 1496 99 1504 102
rect 1431 92 1433 94
rect 1435 92 1438 94
rect 1431 90 1438 92
rect 1499 96 1504 99
rect 1506 96 1511 108
rect 1513 96 1521 108
rect 1525 107 1532 109
rect 1527 104 1532 107
rect 1534 107 1542 113
rect 1544 111 1552 113
rect 1544 109 1547 111
rect 1549 109 1552 111
rect 1544 107 1552 109
rect 1554 107 1561 113
rect 1606 111 1613 113
rect 1567 108 1572 111
rect 1534 104 1540 107
rect 1536 100 1540 104
rect 1556 100 1561 107
rect 1565 106 1572 108
rect 1565 104 1567 106
rect 1569 104 1572 106
rect 1565 102 1572 104
rect 1574 102 1585 111
rect 1536 98 1542 100
rect 1536 96 1538 98
rect 1540 96 1542 98
rect 1515 94 1521 96
rect 1515 92 1517 94
rect 1519 92 1521 94
rect 1515 90 1521 92
rect 1536 94 1542 96
rect 1555 98 1561 100
rect 1576 100 1585 102
rect 1587 100 1592 111
rect 1594 106 1599 111
rect 1606 109 1608 111
rect 1610 109 1613 111
rect 1606 107 1613 109
rect 1594 104 1601 106
rect 1608 104 1613 107
rect 1615 108 1620 113
rect 1711 111 1718 113
rect 1672 108 1677 111
rect 1615 104 1629 108
rect 1594 102 1597 104
rect 1599 102 1601 104
rect 1594 100 1601 102
rect 1620 103 1629 104
rect 1620 101 1622 103
rect 1624 101 1629 103
rect 1555 96 1557 98
rect 1559 96 1561 98
rect 1555 94 1561 96
rect 1576 94 1583 100
rect 1620 99 1629 101
rect 1631 106 1639 108
rect 1631 104 1634 106
rect 1636 104 1639 106
rect 1631 99 1639 104
rect 1641 104 1649 108
rect 1641 102 1644 104
rect 1646 102 1649 104
rect 1641 99 1649 102
rect 1576 92 1578 94
rect 1580 92 1583 94
rect 1576 90 1583 92
rect 1644 96 1649 99
rect 1651 96 1656 108
rect 1658 96 1666 108
rect 1670 106 1677 108
rect 1670 104 1672 106
rect 1674 104 1677 106
rect 1670 102 1677 104
rect 1679 102 1690 111
rect 1681 100 1690 102
rect 1692 100 1697 111
rect 1699 106 1704 111
rect 1711 109 1713 111
rect 1715 109 1718 111
rect 1711 107 1718 109
rect 1699 104 1706 106
rect 1713 104 1718 107
rect 1720 108 1725 113
rect 1944 111 1951 113
rect 1825 108 1830 111
rect 1720 104 1734 108
rect 1699 102 1702 104
rect 1704 102 1706 104
rect 1699 100 1706 102
rect 1725 103 1734 104
rect 1725 101 1727 103
rect 1729 101 1734 103
rect 1660 94 1666 96
rect 1660 92 1662 94
rect 1664 92 1666 94
rect 1660 90 1666 92
rect 1681 94 1688 100
rect 1725 99 1734 101
rect 1736 106 1744 108
rect 1736 104 1739 106
rect 1741 104 1744 106
rect 1736 99 1744 104
rect 1746 104 1754 108
rect 1746 102 1749 104
rect 1751 102 1754 104
rect 1746 99 1754 102
rect 1681 92 1683 94
rect 1685 92 1688 94
rect 1681 90 1688 92
rect 1749 96 1754 99
rect 1756 96 1761 108
rect 1763 96 1771 108
rect 1823 106 1830 108
rect 1823 104 1825 106
rect 1827 104 1830 106
rect 1823 102 1830 104
rect 1832 102 1843 111
rect 1834 100 1843 102
rect 1845 100 1850 111
rect 1852 106 1857 111
rect 1865 106 1870 111
rect 1852 104 1859 106
rect 1852 102 1855 104
rect 1857 102 1859 104
rect 1852 100 1859 102
rect 1863 104 1870 106
rect 1863 102 1865 104
rect 1867 102 1870 104
rect 1863 100 1870 102
rect 1872 100 1877 111
rect 1879 102 1890 111
rect 1892 108 1897 111
rect 1905 108 1910 111
rect 1892 106 1899 108
rect 1892 104 1895 106
rect 1897 104 1899 106
rect 1892 102 1899 104
rect 1903 106 1910 108
rect 1903 104 1905 106
rect 1907 104 1910 106
rect 1903 102 1910 104
rect 1912 102 1923 111
rect 1879 100 1888 102
rect 1765 94 1771 96
rect 1765 92 1767 94
rect 1769 92 1771 94
rect 1765 90 1771 92
rect 1834 94 1841 100
rect 1834 92 1836 94
rect 1838 92 1841 94
rect 1834 90 1841 92
rect 1881 94 1888 100
rect 1914 100 1923 102
rect 1925 100 1930 111
rect 1932 106 1937 111
rect 1944 109 1946 111
rect 1948 109 1951 111
rect 1944 107 1951 109
rect 1932 104 1939 106
rect 1946 104 1951 107
rect 1953 108 1958 113
rect 1953 104 1967 108
rect 1932 102 1935 104
rect 1937 102 1939 104
rect 1932 100 1939 102
rect 1958 103 1967 104
rect 1958 101 1960 103
rect 1962 101 1967 103
rect 1881 92 1884 94
rect 1886 92 1888 94
rect 1881 90 1888 92
rect 1914 94 1921 100
rect 1958 99 1967 101
rect 1969 106 1977 108
rect 1969 104 1972 106
rect 1974 104 1977 106
rect 1969 99 1977 104
rect 1979 104 1987 108
rect 1979 102 1982 104
rect 1984 102 1987 104
rect 1979 99 1987 102
rect 1914 92 1916 94
rect 1918 92 1921 94
rect 1914 90 1921 92
rect 1982 96 1987 99
rect 1989 96 1994 108
rect 1996 96 2004 108
rect 1998 94 2004 96
rect 1998 92 2000 94
rect 2002 92 2004 94
rect 1998 90 2004 92
rect 18 68 24 70
rect 18 66 20 68
rect 22 66 24 68
rect 18 64 24 66
rect 37 68 43 70
rect 58 72 65 74
rect 58 70 60 72
rect 62 70 65 72
rect 37 66 39 68
rect 41 66 43 68
rect 37 64 43 66
rect 18 60 22 64
rect 9 57 14 60
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect 7 51 14 53
rect 16 57 22 60
rect 38 57 43 64
rect 58 64 65 70
rect 142 72 148 74
rect 142 70 144 72
rect 146 70 148 72
rect 142 68 148 70
rect 163 72 170 74
rect 163 70 165 72
rect 167 70 170 72
rect 126 65 131 68
rect 58 62 67 64
rect 16 51 24 57
rect 26 55 34 57
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 51 43 57
rect 47 60 54 62
rect 47 58 49 60
rect 51 58 54 60
rect 47 56 54 58
rect 49 53 54 56
rect 56 53 67 62
rect 69 53 74 64
rect 76 62 83 64
rect 76 60 79 62
rect 81 60 83 62
rect 102 63 111 65
rect 102 61 104 63
rect 106 61 111 63
rect 102 60 111 61
rect 76 58 83 60
rect 76 53 81 58
rect 90 57 95 60
rect 88 55 95 57
rect 88 53 90 55
rect 92 53 95 55
rect 88 51 95 53
rect 97 56 111 60
rect 113 60 121 65
rect 113 58 116 60
rect 118 58 121 60
rect 113 56 121 58
rect 123 62 131 65
rect 123 60 126 62
rect 128 60 131 62
rect 123 56 131 60
rect 133 56 138 68
rect 140 56 148 68
rect 163 64 170 70
rect 247 72 253 74
rect 247 70 249 72
rect 251 70 253 72
rect 247 68 253 70
rect 268 68 274 70
rect 231 65 236 68
rect 163 62 172 64
rect 152 60 159 62
rect 152 58 154 60
rect 156 58 159 60
rect 152 56 159 58
rect 97 51 102 56
rect 154 53 159 56
rect 161 53 172 62
rect 174 53 179 64
rect 181 62 188 64
rect 181 60 184 62
rect 186 60 188 62
rect 207 63 216 65
rect 207 61 209 63
rect 211 61 216 63
rect 207 60 216 61
rect 181 58 188 60
rect 181 53 186 58
rect 195 57 200 60
rect 193 55 200 57
rect 193 53 195 55
rect 197 53 200 55
rect 193 51 200 53
rect 202 56 216 60
rect 218 60 226 65
rect 218 58 221 60
rect 223 58 226 60
rect 218 56 226 58
rect 228 62 236 65
rect 228 60 231 62
rect 233 60 236 62
rect 228 56 236 60
rect 238 56 243 68
rect 245 56 253 68
rect 268 66 270 68
rect 272 66 274 68
rect 268 64 274 66
rect 287 68 293 70
rect 308 72 315 74
rect 308 70 310 72
rect 312 70 315 72
rect 287 66 289 68
rect 291 66 293 68
rect 287 64 293 66
rect 268 60 272 64
rect 259 57 264 60
rect 202 51 207 56
rect 257 55 264 57
rect 257 53 259 55
rect 261 53 264 55
rect 257 51 264 53
rect 266 57 272 60
rect 288 57 293 64
rect 308 64 315 70
rect 392 72 398 74
rect 392 70 394 72
rect 396 70 398 72
rect 392 68 398 70
rect 413 72 420 74
rect 413 70 415 72
rect 417 70 420 72
rect 376 65 381 68
rect 308 62 317 64
rect 266 51 274 57
rect 276 55 284 57
rect 276 53 279 55
rect 281 53 284 55
rect 276 51 284 53
rect 286 51 293 57
rect 297 60 304 62
rect 297 58 299 60
rect 301 58 304 60
rect 297 56 304 58
rect 299 53 304 56
rect 306 53 317 62
rect 319 53 324 64
rect 326 62 333 64
rect 326 60 329 62
rect 331 60 333 62
rect 352 63 361 65
rect 352 61 354 63
rect 356 61 361 63
rect 352 60 361 61
rect 326 58 333 60
rect 326 53 331 58
rect 340 57 345 60
rect 338 55 345 57
rect 338 53 340 55
rect 342 53 345 55
rect 338 51 345 53
rect 347 56 361 60
rect 363 60 371 65
rect 363 58 366 60
rect 368 58 371 60
rect 363 56 371 58
rect 373 62 381 65
rect 373 60 376 62
rect 378 60 381 62
rect 373 56 381 60
rect 383 56 388 68
rect 390 56 398 68
rect 413 64 420 70
rect 497 72 503 74
rect 497 70 499 72
rect 501 70 503 72
rect 497 68 503 70
rect 518 68 524 70
rect 481 65 486 68
rect 413 62 422 64
rect 402 60 409 62
rect 402 58 404 60
rect 406 58 409 60
rect 402 56 409 58
rect 347 51 352 56
rect 404 53 409 56
rect 411 53 422 62
rect 424 53 429 64
rect 431 62 438 64
rect 431 60 434 62
rect 436 60 438 62
rect 457 63 466 65
rect 457 61 459 63
rect 461 61 466 63
rect 457 60 466 61
rect 431 58 438 60
rect 431 53 436 58
rect 445 57 450 60
rect 443 55 450 57
rect 443 53 445 55
rect 447 53 450 55
rect 443 51 450 53
rect 452 56 466 60
rect 468 60 476 65
rect 468 58 471 60
rect 473 58 476 60
rect 468 56 476 58
rect 478 62 486 65
rect 478 60 481 62
rect 483 60 486 62
rect 478 56 486 60
rect 488 56 493 68
rect 495 56 503 68
rect 518 66 520 68
rect 522 66 524 68
rect 518 64 524 66
rect 537 68 543 70
rect 558 72 565 74
rect 558 70 560 72
rect 562 70 565 72
rect 537 66 539 68
rect 541 66 543 68
rect 537 64 543 66
rect 518 60 522 64
rect 509 57 514 60
rect 452 51 457 56
rect 507 55 514 57
rect 507 53 509 55
rect 511 53 514 55
rect 507 51 514 53
rect 516 57 522 60
rect 538 57 543 64
rect 558 64 565 70
rect 642 72 648 74
rect 642 70 644 72
rect 646 70 648 72
rect 642 68 648 70
rect 663 72 670 74
rect 663 70 665 72
rect 667 70 670 72
rect 626 65 631 68
rect 558 62 567 64
rect 516 51 524 57
rect 526 55 534 57
rect 526 53 529 55
rect 531 53 534 55
rect 526 51 534 53
rect 536 51 543 57
rect 547 60 554 62
rect 547 58 549 60
rect 551 58 554 60
rect 547 56 554 58
rect 549 53 554 56
rect 556 53 567 62
rect 569 53 574 64
rect 576 62 583 64
rect 576 60 579 62
rect 581 60 583 62
rect 602 63 611 65
rect 602 61 604 63
rect 606 61 611 63
rect 602 60 611 61
rect 576 58 583 60
rect 576 53 581 58
rect 590 57 595 60
rect 588 55 595 57
rect 588 53 590 55
rect 592 53 595 55
rect 588 51 595 53
rect 597 56 611 60
rect 613 60 621 65
rect 613 58 616 60
rect 618 58 621 60
rect 613 56 621 58
rect 623 62 631 65
rect 623 60 626 62
rect 628 60 631 62
rect 623 56 631 60
rect 633 56 638 68
rect 640 56 648 68
rect 663 64 670 70
rect 747 72 753 74
rect 747 70 749 72
rect 751 70 753 72
rect 747 68 753 70
rect 768 68 774 70
rect 731 65 736 68
rect 663 62 672 64
rect 652 60 659 62
rect 652 58 654 60
rect 656 58 659 60
rect 652 56 659 58
rect 597 51 602 56
rect 654 53 659 56
rect 661 53 672 62
rect 674 53 679 64
rect 681 62 688 64
rect 681 60 684 62
rect 686 60 688 62
rect 707 63 716 65
rect 707 61 709 63
rect 711 61 716 63
rect 707 60 716 61
rect 681 58 688 60
rect 681 53 686 58
rect 695 57 700 60
rect 693 55 700 57
rect 693 53 695 55
rect 697 53 700 55
rect 693 51 700 53
rect 702 56 716 60
rect 718 60 726 65
rect 718 58 721 60
rect 723 58 726 60
rect 718 56 726 58
rect 728 62 736 65
rect 728 60 731 62
rect 733 60 736 62
rect 728 56 736 60
rect 738 56 743 68
rect 745 56 753 68
rect 768 66 770 68
rect 772 66 774 68
rect 768 64 774 66
rect 787 68 793 70
rect 808 72 815 74
rect 808 70 810 72
rect 812 70 815 72
rect 787 66 789 68
rect 791 66 793 68
rect 787 64 793 66
rect 768 60 772 64
rect 759 57 764 60
rect 702 51 707 56
rect 757 55 764 57
rect 757 53 759 55
rect 761 53 764 55
rect 757 51 764 53
rect 766 57 772 60
rect 788 57 793 64
rect 808 64 815 70
rect 892 72 898 74
rect 892 70 894 72
rect 896 70 898 72
rect 892 68 898 70
rect 913 72 920 74
rect 913 70 915 72
rect 917 70 920 72
rect 876 65 881 68
rect 808 62 817 64
rect 766 51 774 57
rect 776 55 784 57
rect 776 53 779 55
rect 781 53 784 55
rect 776 51 784 53
rect 786 51 793 57
rect 797 60 804 62
rect 797 58 799 60
rect 801 58 804 60
rect 797 56 804 58
rect 799 53 804 56
rect 806 53 817 62
rect 819 53 824 64
rect 826 62 833 64
rect 826 60 829 62
rect 831 60 833 62
rect 852 63 861 65
rect 852 61 854 63
rect 856 61 861 63
rect 852 60 861 61
rect 826 58 833 60
rect 826 53 831 58
rect 840 57 845 60
rect 838 55 845 57
rect 838 53 840 55
rect 842 53 845 55
rect 838 51 845 53
rect 847 56 861 60
rect 863 60 871 65
rect 863 58 866 60
rect 868 58 871 60
rect 863 56 871 58
rect 873 62 881 65
rect 873 60 876 62
rect 878 60 881 62
rect 873 56 881 60
rect 883 56 888 68
rect 890 56 898 68
rect 913 64 920 70
rect 997 72 1003 74
rect 997 70 999 72
rect 1001 70 1003 72
rect 997 68 1003 70
rect 1028 68 1034 70
rect 981 65 986 68
rect 913 62 922 64
rect 902 60 909 62
rect 902 58 904 60
rect 906 58 909 60
rect 902 56 909 58
rect 847 51 852 56
rect 904 53 909 56
rect 911 53 922 62
rect 924 53 929 64
rect 931 62 938 64
rect 931 60 934 62
rect 936 60 938 62
rect 957 63 966 65
rect 957 61 959 63
rect 961 61 966 63
rect 957 60 966 61
rect 931 58 938 60
rect 931 53 936 58
rect 945 57 950 60
rect 943 55 950 57
rect 943 53 945 55
rect 947 53 950 55
rect 943 51 950 53
rect 952 56 966 60
rect 968 60 976 65
rect 968 58 971 60
rect 973 58 976 60
rect 968 56 976 58
rect 978 62 986 65
rect 978 60 981 62
rect 983 60 986 62
rect 978 56 986 60
rect 988 56 993 68
rect 995 56 1003 68
rect 1028 66 1030 68
rect 1032 66 1034 68
rect 1028 64 1034 66
rect 1047 68 1053 70
rect 1068 72 1075 74
rect 1068 70 1070 72
rect 1072 70 1075 72
rect 1047 66 1049 68
rect 1051 66 1053 68
rect 1047 64 1053 66
rect 1028 60 1032 64
rect 1019 57 1024 60
rect 952 51 957 56
rect 1017 55 1024 57
rect 1017 53 1019 55
rect 1021 53 1024 55
rect 1017 51 1024 53
rect 1026 57 1032 60
rect 1048 57 1053 64
rect 1068 64 1075 70
rect 1152 72 1158 74
rect 1152 70 1154 72
rect 1156 70 1158 72
rect 1152 68 1158 70
rect 1173 72 1180 74
rect 1173 70 1175 72
rect 1177 70 1180 72
rect 1136 65 1141 68
rect 1068 62 1077 64
rect 1026 51 1034 57
rect 1036 55 1044 57
rect 1036 53 1039 55
rect 1041 53 1044 55
rect 1036 51 1044 53
rect 1046 51 1053 57
rect 1057 60 1064 62
rect 1057 58 1059 60
rect 1061 58 1064 60
rect 1057 56 1064 58
rect 1059 53 1064 56
rect 1066 53 1077 62
rect 1079 53 1084 64
rect 1086 62 1093 64
rect 1086 60 1089 62
rect 1091 60 1093 62
rect 1112 63 1121 65
rect 1112 61 1114 63
rect 1116 61 1121 63
rect 1112 60 1121 61
rect 1086 58 1093 60
rect 1086 53 1091 58
rect 1100 57 1105 60
rect 1098 55 1105 57
rect 1098 53 1100 55
rect 1102 53 1105 55
rect 1098 51 1105 53
rect 1107 56 1121 60
rect 1123 60 1131 65
rect 1123 58 1126 60
rect 1128 58 1131 60
rect 1123 56 1131 58
rect 1133 62 1141 65
rect 1133 60 1136 62
rect 1138 60 1141 62
rect 1133 56 1141 60
rect 1143 56 1148 68
rect 1150 56 1158 68
rect 1173 64 1180 70
rect 1257 72 1263 74
rect 1257 70 1259 72
rect 1261 70 1263 72
rect 1257 68 1263 70
rect 1278 68 1284 70
rect 1241 65 1246 68
rect 1173 62 1182 64
rect 1162 60 1169 62
rect 1162 58 1164 60
rect 1166 58 1169 60
rect 1162 56 1169 58
rect 1107 51 1112 56
rect 1164 53 1169 56
rect 1171 53 1182 62
rect 1184 53 1189 64
rect 1191 62 1198 64
rect 1191 60 1194 62
rect 1196 60 1198 62
rect 1217 63 1226 65
rect 1217 61 1219 63
rect 1221 61 1226 63
rect 1217 60 1226 61
rect 1191 58 1198 60
rect 1191 53 1196 58
rect 1205 57 1210 60
rect 1203 55 1210 57
rect 1203 53 1205 55
rect 1207 53 1210 55
rect 1203 51 1210 53
rect 1212 56 1226 60
rect 1228 60 1236 65
rect 1228 58 1231 60
rect 1233 58 1236 60
rect 1228 56 1236 58
rect 1238 62 1246 65
rect 1238 60 1241 62
rect 1243 60 1246 62
rect 1238 56 1246 60
rect 1248 56 1253 68
rect 1255 56 1263 68
rect 1278 66 1280 68
rect 1282 66 1284 68
rect 1278 64 1284 66
rect 1297 68 1303 70
rect 1318 72 1325 74
rect 1318 70 1320 72
rect 1322 70 1325 72
rect 1297 66 1299 68
rect 1301 66 1303 68
rect 1297 64 1303 66
rect 1278 60 1282 64
rect 1269 57 1274 60
rect 1212 51 1217 56
rect 1267 55 1274 57
rect 1267 53 1269 55
rect 1271 53 1274 55
rect 1267 51 1274 53
rect 1276 57 1282 60
rect 1298 57 1303 64
rect 1318 64 1325 70
rect 1402 72 1408 74
rect 1402 70 1404 72
rect 1406 70 1408 72
rect 1402 68 1408 70
rect 1423 72 1430 74
rect 1423 70 1425 72
rect 1427 70 1430 72
rect 1386 65 1391 68
rect 1318 62 1327 64
rect 1276 51 1284 57
rect 1286 55 1294 57
rect 1286 53 1289 55
rect 1291 53 1294 55
rect 1286 51 1294 53
rect 1296 51 1303 57
rect 1307 60 1314 62
rect 1307 58 1309 60
rect 1311 58 1314 60
rect 1307 56 1314 58
rect 1309 53 1314 56
rect 1316 53 1327 62
rect 1329 53 1334 64
rect 1336 62 1343 64
rect 1336 60 1339 62
rect 1341 60 1343 62
rect 1362 63 1371 65
rect 1362 61 1364 63
rect 1366 61 1371 63
rect 1362 60 1371 61
rect 1336 58 1343 60
rect 1336 53 1341 58
rect 1350 57 1355 60
rect 1348 55 1355 57
rect 1348 53 1350 55
rect 1352 53 1355 55
rect 1348 51 1355 53
rect 1357 56 1371 60
rect 1373 60 1381 65
rect 1373 58 1376 60
rect 1378 58 1381 60
rect 1373 56 1381 58
rect 1383 62 1391 65
rect 1383 60 1386 62
rect 1388 60 1391 62
rect 1383 56 1391 60
rect 1393 56 1398 68
rect 1400 56 1408 68
rect 1423 64 1430 70
rect 1507 72 1513 74
rect 1507 70 1509 72
rect 1511 70 1513 72
rect 1507 68 1513 70
rect 1528 68 1534 70
rect 1491 65 1496 68
rect 1423 62 1432 64
rect 1412 60 1419 62
rect 1412 58 1414 60
rect 1416 58 1419 60
rect 1412 56 1419 58
rect 1357 51 1362 56
rect 1414 53 1419 56
rect 1421 53 1432 62
rect 1434 53 1439 64
rect 1441 62 1448 64
rect 1441 60 1444 62
rect 1446 60 1448 62
rect 1467 63 1476 65
rect 1467 61 1469 63
rect 1471 61 1476 63
rect 1467 60 1476 61
rect 1441 58 1448 60
rect 1441 53 1446 58
rect 1455 57 1460 60
rect 1453 55 1460 57
rect 1453 53 1455 55
rect 1457 53 1460 55
rect 1453 51 1460 53
rect 1462 56 1476 60
rect 1478 60 1486 65
rect 1478 58 1481 60
rect 1483 58 1486 60
rect 1478 56 1486 58
rect 1488 62 1496 65
rect 1488 60 1491 62
rect 1493 60 1496 62
rect 1488 56 1496 60
rect 1498 56 1503 68
rect 1505 56 1513 68
rect 1528 66 1530 68
rect 1532 66 1534 68
rect 1528 64 1534 66
rect 1547 68 1553 70
rect 1568 72 1575 74
rect 1568 70 1570 72
rect 1572 70 1575 72
rect 1547 66 1549 68
rect 1551 66 1553 68
rect 1547 64 1553 66
rect 1528 60 1532 64
rect 1519 57 1524 60
rect 1462 51 1467 56
rect 1517 55 1524 57
rect 1517 53 1519 55
rect 1521 53 1524 55
rect 1517 51 1524 53
rect 1526 57 1532 60
rect 1548 57 1553 64
rect 1568 64 1575 70
rect 1652 72 1658 74
rect 1652 70 1654 72
rect 1656 70 1658 72
rect 1652 68 1658 70
rect 1673 72 1680 74
rect 1673 70 1675 72
rect 1677 70 1680 72
rect 1636 65 1641 68
rect 1568 62 1577 64
rect 1526 51 1534 57
rect 1536 55 1544 57
rect 1536 53 1539 55
rect 1541 53 1544 55
rect 1536 51 1544 53
rect 1546 51 1553 57
rect 1557 60 1564 62
rect 1557 58 1559 60
rect 1561 58 1564 60
rect 1557 56 1564 58
rect 1559 53 1564 56
rect 1566 53 1577 62
rect 1579 53 1584 64
rect 1586 62 1593 64
rect 1586 60 1589 62
rect 1591 60 1593 62
rect 1612 63 1621 65
rect 1612 61 1614 63
rect 1616 61 1621 63
rect 1612 60 1621 61
rect 1586 58 1593 60
rect 1586 53 1591 58
rect 1600 57 1605 60
rect 1598 55 1605 57
rect 1598 53 1600 55
rect 1602 53 1605 55
rect 1598 51 1605 53
rect 1607 56 1621 60
rect 1623 60 1631 65
rect 1623 58 1626 60
rect 1628 58 1631 60
rect 1623 56 1631 58
rect 1633 62 1641 65
rect 1633 60 1636 62
rect 1638 60 1641 62
rect 1633 56 1641 60
rect 1643 56 1648 68
rect 1650 56 1658 68
rect 1673 64 1680 70
rect 1757 72 1763 74
rect 1757 70 1759 72
rect 1761 70 1763 72
rect 1757 68 1763 70
rect 1778 68 1784 70
rect 1741 65 1746 68
rect 1673 62 1682 64
rect 1662 60 1669 62
rect 1662 58 1664 60
rect 1666 58 1669 60
rect 1662 56 1669 58
rect 1607 51 1612 56
rect 1664 53 1669 56
rect 1671 53 1682 62
rect 1684 53 1689 64
rect 1691 62 1698 64
rect 1691 60 1694 62
rect 1696 60 1698 62
rect 1717 63 1726 65
rect 1717 61 1719 63
rect 1721 61 1726 63
rect 1717 60 1726 61
rect 1691 58 1698 60
rect 1691 53 1696 58
rect 1705 57 1710 60
rect 1703 55 1710 57
rect 1703 53 1705 55
rect 1707 53 1710 55
rect 1703 51 1710 53
rect 1712 56 1726 60
rect 1728 60 1736 65
rect 1728 58 1731 60
rect 1733 58 1736 60
rect 1728 56 1736 58
rect 1738 62 1746 65
rect 1738 60 1741 62
rect 1743 60 1746 62
rect 1738 56 1746 60
rect 1748 56 1753 68
rect 1755 56 1763 68
rect 1778 66 1780 68
rect 1782 66 1784 68
rect 1778 64 1784 66
rect 1797 68 1803 70
rect 1818 72 1825 74
rect 1818 70 1820 72
rect 1822 70 1825 72
rect 1797 66 1799 68
rect 1801 66 1803 68
rect 1797 64 1803 66
rect 1778 60 1782 64
rect 1769 57 1774 60
rect 1712 51 1717 56
rect 1767 55 1774 57
rect 1767 53 1769 55
rect 1771 53 1774 55
rect 1767 51 1774 53
rect 1776 57 1782 60
rect 1798 57 1803 64
rect 1818 64 1825 70
rect 1902 72 1908 74
rect 1902 70 1904 72
rect 1906 70 1908 72
rect 1902 68 1908 70
rect 1923 72 1930 74
rect 1923 70 1925 72
rect 1927 70 1930 72
rect 1886 65 1891 68
rect 1818 62 1827 64
rect 1776 51 1784 57
rect 1786 55 1794 57
rect 1786 53 1789 55
rect 1791 53 1794 55
rect 1786 51 1794 53
rect 1796 51 1803 57
rect 1807 60 1814 62
rect 1807 58 1809 60
rect 1811 58 1814 60
rect 1807 56 1814 58
rect 1809 53 1814 56
rect 1816 53 1827 62
rect 1829 53 1834 64
rect 1836 62 1843 64
rect 1836 60 1839 62
rect 1841 60 1843 62
rect 1862 63 1871 65
rect 1862 61 1864 63
rect 1866 61 1871 63
rect 1862 60 1871 61
rect 1836 58 1843 60
rect 1836 53 1841 58
rect 1850 57 1855 60
rect 1848 55 1855 57
rect 1848 53 1850 55
rect 1852 53 1855 55
rect 1848 51 1855 53
rect 1857 56 1871 60
rect 1873 60 1881 65
rect 1873 58 1876 60
rect 1878 58 1881 60
rect 1873 56 1881 58
rect 1883 62 1891 65
rect 1883 60 1886 62
rect 1888 60 1891 62
rect 1883 56 1891 60
rect 1893 56 1898 68
rect 1900 56 1908 68
rect 1923 64 1930 70
rect 2007 72 2013 74
rect 2007 70 2009 72
rect 2011 70 2013 72
rect 2007 68 2013 70
rect 1991 65 1996 68
rect 1923 62 1932 64
rect 1912 60 1919 62
rect 1912 58 1914 60
rect 1916 58 1919 60
rect 1912 56 1919 58
rect 1857 51 1862 56
rect 1914 53 1919 56
rect 1921 53 1932 62
rect 1934 53 1939 64
rect 1941 62 1948 64
rect 1941 60 1944 62
rect 1946 60 1948 62
rect 1967 63 1976 65
rect 1967 61 1969 63
rect 1971 61 1976 63
rect 1967 60 1976 61
rect 1941 58 1948 60
rect 1941 53 1946 58
rect 1955 57 1960 60
rect 1953 55 1960 57
rect 1953 53 1955 55
rect 1957 53 1960 55
rect 1953 51 1960 53
rect 1962 56 1976 60
rect 1978 60 1986 65
rect 1978 58 1981 60
rect 1983 58 1986 60
rect 1978 56 1986 58
rect 1988 62 1996 65
rect 1988 60 1991 62
rect 1993 60 1996 62
rect 1988 56 1996 60
rect 1998 56 2003 68
rect 2005 56 2013 68
rect 1962 51 1967 56
<< pdif >>
rect 54 185 60 192
rect 33 176 40 185
rect 33 174 35 176
rect 37 174 40 176
rect 33 172 40 174
rect 42 183 50 185
rect 42 181 45 183
rect 47 181 50 183
rect 42 176 50 181
rect 42 174 45 176
rect 47 174 50 176
rect 42 172 50 174
rect 52 178 60 185
rect 52 176 55 178
rect 57 176 60 178
rect 52 174 60 176
rect 62 190 69 192
rect 62 188 65 190
rect 67 188 69 190
rect 62 183 69 188
rect 94 185 100 192
rect 62 181 65 183
rect 67 181 69 183
rect 62 179 69 181
rect 62 174 67 179
rect 73 176 80 185
rect 73 174 75 176
rect 77 174 80 176
rect 52 172 58 174
rect 73 172 80 174
rect 82 183 90 185
rect 82 181 85 183
rect 87 181 90 183
rect 82 176 90 181
rect 82 174 85 176
rect 87 174 90 176
rect 82 172 90 174
rect 92 178 100 185
rect 92 176 95 178
rect 97 176 100 178
rect 92 174 100 176
rect 102 190 109 192
rect 102 188 105 190
rect 107 188 109 190
rect 102 183 109 188
rect 102 181 105 183
rect 107 181 109 183
rect 102 179 109 181
rect 102 174 107 179
rect 122 177 127 192
rect 120 175 127 177
rect 92 172 98 174
rect 120 173 122 175
rect 124 173 127 175
rect 120 171 127 173
rect 122 165 127 171
rect 129 183 137 192
rect 129 181 132 183
rect 134 181 137 183
rect 129 174 137 181
rect 139 190 147 192
rect 139 188 142 190
rect 144 188 147 190
rect 139 183 147 188
rect 139 181 142 183
rect 144 181 147 183
rect 139 174 147 181
rect 149 176 163 192
rect 149 174 158 176
rect 160 174 163 176
rect 129 165 134 174
rect 151 169 163 174
rect 151 167 158 169
rect 160 167 163 169
rect 151 165 163 167
rect 165 190 172 192
rect 165 188 168 190
rect 170 188 172 190
rect 165 186 172 188
rect 165 165 170 186
rect 206 185 212 192
rect 185 176 192 185
rect 185 174 187 176
rect 189 174 192 176
rect 185 172 192 174
rect 194 183 202 185
rect 194 181 197 183
rect 199 181 202 183
rect 194 176 202 181
rect 194 174 197 176
rect 199 174 202 176
rect 194 172 202 174
rect 204 178 212 185
rect 204 176 207 178
rect 209 176 212 178
rect 204 174 212 176
rect 214 190 221 192
rect 214 188 217 190
rect 219 188 221 190
rect 214 183 221 188
rect 214 181 217 183
rect 219 181 221 183
rect 214 179 221 181
rect 363 189 370 191
rect 363 187 365 189
rect 367 187 370 189
rect 363 182 370 187
rect 363 180 365 182
rect 367 180 370 182
rect 214 174 219 179
rect 363 178 370 180
rect 204 172 210 174
rect 365 173 370 178
rect 372 184 378 191
rect 424 184 430 191
rect 372 177 380 184
rect 372 175 375 177
rect 377 175 380 177
rect 372 173 380 175
rect 374 171 380 173
rect 382 182 390 184
rect 382 180 385 182
rect 387 180 390 182
rect 382 175 390 180
rect 382 173 385 175
rect 387 173 390 175
rect 382 171 390 173
rect 392 175 399 184
rect 392 173 395 175
rect 397 173 399 175
rect 392 171 399 173
rect 403 175 410 184
rect 403 173 405 175
rect 407 173 410 175
rect 403 171 410 173
rect 412 182 420 184
rect 412 180 415 182
rect 417 180 420 182
rect 412 175 420 180
rect 412 173 415 175
rect 417 173 420 175
rect 412 171 420 173
rect 422 177 430 184
rect 422 175 425 177
rect 427 175 430 177
rect 422 173 430 175
rect 432 189 439 191
rect 432 187 435 189
rect 437 187 439 189
rect 432 182 439 187
rect 432 180 435 182
rect 437 180 439 182
rect 432 178 439 180
rect 443 189 450 191
rect 443 187 445 189
rect 447 187 450 189
rect 443 182 450 187
rect 443 180 445 182
rect 447 180 450 182
rect 443 178 450 180
rect 432 173 437 178
rect 445 173 450 178
rect 452 184 458 191
rect 492 189 499 191
rect 492 187 494 189
rect 496 187 499 189
rect 492 185 499 187
rect 452 177 460 184
rect 452 175 455 177
rect 457 175 460 177
rect 452 173 460 175
rect 422 171 428 173
rect 454 171 460 173
rect 462 182 470 184
rect 462 180 465 182
rect 467 180 470 182
rect 462 175 470 180
rect 462 173 465 175
rect 467 173 470 175
rect 462 171 470 173
rect 472 175 479 184
rect 472 173 475 175
rect 477 173 479 175
rect 472 171 479 173
rect 494 164 499 185
rect 501 175 515 191
rect 501 173 504 175
rect 506 173 515 175
rect 517 189 525 191
rect 517 187 520 189
rect 522 187 525 189
rect 517 182 525 187
rect 517 180 520 182
rect 522 180 525 182
rect 517 173 525 180
rect 527 182 535 191
rect 527 180 530 182
rect 532 180 535 182
rect 527 173 535 180
rect 501 168 513 173
rect 501 166 504 168
rect 506 166 513 168
rect 501 164 513 166
rect 530 164 535 173
rect 537 176 542 191
rect 568 189 575 191
rect 568 187 570 189
rect 572 187 575 189
rect 568 182 575 187
rect 568 180 570 182
rect 572 180 575 182
rect 568 178 575 180
rect 537 174 544 176
rect 537 172 540 174
rect 542 172 544 174
rect 570 173 575 178
rect 577 184 583 191
rect 629 184 635 191
rect 577 177 585 184
rect 577 175 580 177
rect 582 175 585 177
rect 577 173 585 175
rect 537 170 544 172
rect 537 164 542 170
rect 579 171 585 173
rect 587 182 595 184
rect 587 180 590 182
rect 592 180 595 182
rect 587 175 595 180
rect 587 173 590 175
rect 592 173 595 175
rect 587 171 595 173
rect 597 175 604 184
rect 597 173 600 175
rect 602 173 604 175
rect 597 171 604 173
rect 608 175 615 184
rect 608 173 610 175
rect 612 173 615 175
rect 608 171 615 173
rect 617 182 625 184
rect 617 180 620 182
rect 622 180 625 182
rect 617 175 625 180
rect 617 173 620 175
rect 622 173 625 175
rect 617 171 625 173
rect 627 177 635 184
rect 627 175 630 177
rect 632 175 635 177
rect 627 173 635 175
rect 637 189 644 191
rect 637 187 640 189
rect 642 187 644 189
rect 637 182 644 187
rect 637 180 640 182
rect 642 180 644 182
rect 637 178 644 180
rect 648 189 655 191
rect 648 187 650 189
rect 652 187 655 189
rect 648 182 655 187
rect 648 180 650 182
rect 652 180 655 182
rect 648 178 655 180
rect 637 173 642 178
rect 650 173 655 178
rect 657 184 663 191
rect 697 189 704 191
rect 697 187 699 189
rect 701 187 704 189
rect 697 185 704 187
rect 657 177 665 184
rect 657 175 660 177
rect 662 175 665 177
rect 657 173 665 175
rect 627 171 633 173
rect 659 171 665 173
rect 667 182 675 184
rect 667 180 670 182
rect 672 180 675 182
rect 667 175 675 180
rect 667 173 670 175
rect 672 173 675 175
rect 667 171 675 173
rect 677 175 684 184
rect 677 173 680 175
rect 682 173 684 175
rect 677 171 684 173
rect 699 164 704 185
rect 706 175 720 191
rect 706 173 709 175
rect 711 173 720 175
rect 722 189 730 191
rect 722 187 725 189
rect 727 187 730 189
rect 722 182 730 187
rect 722 180 725 182
rect 727 180 730 182
rect 722 173 730 180
rect 732 182 740 191
rect 732 180 735 182
rect 737 180 740 182
rect 732 173 740 180
rect 706 168 718 173
rect 706 166 709 168
rect 711 166 718 168
rect 706 164 718 166
rect 735 164 740 173
rect 742 176 747 191
rect 1844 185 1850 192
rect 1823 176 1830 185
rect 742 174 749 176
rect 742 172 745 174
rect 747 172 749 174
rect 1823 174 1825 176
rect 1827 174 1830 176
rect 1823 172 1830 174
rect 1832 183 1840 185
rect 1832 181 1835 183
rect 1837 181 1840 183
rect 1832 176 1840 181
rect 1832 174 1835 176
rect 1837 174 1840 176
rect 1832 172 1840 174
rect 1842 178 1850 185
rect 1842 176 1845 178
rect 1847 176 1850 178
rect 1842 174 1850 176
rect 1852 190 1859 192
rect 1852 188 1855 190
rect 1857 188 1859 190
rect 1852 183 1859 188
rect 1884 185 1890 192
rect 1852 181 1855 183
rect 1857 181 1859 183
rect 1852 179 1859 181
rect 1852 174 1857 179
rect 1863 176 1870 185
rect 1863 174 1865 176
rect 1867 174 1870 176
rect 1842 172 1848 174
rect 742 170 749 172
rect 742 164 747 170
rect 1863 172 1870 174
rect 1872 183 1880 185
rect 1872 181 1875 183
rect 1877 181 1880 183
rect 1872 176 1880 181
rect 1872 174 1875 176
rect 1877 174 1880 176
rect 1872 172 1880 174
rect 1882 178 1890 185
rect 1882 176 1885 178
rect 1887 176 1890 178
rect 1882 174 1890 176
rect 1892 190 1899 192
rect 1892 188 1895 190
rect 1897 188 1899 190
rect 1892 183 1899 188
rect 1892 181 1895 183
rect 1897 181 1899 183
rect 1892 179 1899 181
rect 1892 174 1897 179
rect 1912 177 1917 192
rect 1910 175 1917 177
rect 1882 172 1888 174
rect 1910 173 1912 175
rect 1914 173 1917 175
rect 1910 171 1917 173
rect 1912 165 1917 171
rect 1919 183 1927 192
rect 1919 181 1922 183
rect 1924 181 1927 183
rect 1919 174 1927 181
rect 1929 190 1937 192
rect 1929 188 1932 190
rect 1934 188 1937 190
rect 1929 183 1937 188
rect 1929 181 1932 183
rect 1934 181 1937 183
rect 1929 174 1937 181
rect 1939 176 1953 192
rect 1939 174 1948 176
rect 1950 174 1953 176
rect 1919 165 1924 174
rect 1941 169 1953 174
rect 1941 167 1948 169
rect 1950 167 1953 169
rect 1941 165 1953 167
rect 1955 190 1962 192
rect 1955 188 1958 190
rect 1960 188 1962 190
rect 1955 186 1962 188
rect 1955 165 1960 186
rect 1996 185 2002 192
rect 1975 176 1982 185
rect 1975 174 1977 176
rect 1979 174 1982 176
rect 1975 172 1982 174
rect 1984 183 1992 185
rect 1984 181 1987 183
rect 1989 181 1992 183
rect 1984 176 1992 181
rect 1984 174 1987 176
rect 1989 174 1992 176
rect 1984 172 1992 174
rect 1994 178 2002 185
rect 1994 176 1997 178
rect 1999 176 2002 178
rect 1994 174 2002 176
rect 2004 190 2011 192
rect 2004 188 2007 190
rect 2009 188 2011 190
rect 2004 183 2011 188
rect 2004 181 2007 183
rect 2009 181 2011 183
rect 2004 179 2011 181
rect 2004 174 2009 179
rect 1994 172 2000 174
rect 44 144 50 146
rect 35 139 40 144
rect 33 137 40 139
rect 33 135 35 137
rect 37 135 40 137
rect 33 130 40 135
rect 33 128 35 130
rect 37 128 40 130
rect 33 126 40 128
rect 42 142 50 144
rect 42 140 45 142
rect 47 140 50 142
rect 42 133 50 140
rect 52 144 60 146
rect 52 142 55 144
rect 57 142 60 144
rect 52 137 60 142
rect 52 135 55 137
rect 57 135 60 137
rect 52 133 60 135
rect 62 144 69 146
rect 62 142 65 144
rect 67 142 69 144
rect 62 133 69 142
rect 73 144 80 146
rect 73 142 75 144
rect 77 142 80 144
rect 73 133 80 142
rect 82 144 90 146
rect 82 142 85 144
rect 87 142 90 144
rect 82 137 90 142
rect 82 135 85 137
rect 87 135 90 137
rect 82 133 90 135
rect 92 144 98 146
rect 124 144 130 146
rect 92 142 100 144
rect 92 140 95 142
rect 97 140 100 142
rect 92 133 100 140
rect 42 126 48 133
rect 94 126 100 133
rect 102 139 107 144
rect 115 139 120 144
rect 102 137 109 139
rect 102 135 105 137
rect 107 135 109 137
rect 102 130 109 135
rect 102 128 105 130
rect 107 128 109 130
rect 102 126 109 128
rect 113 137 120 139
rect 113 135 115 137
rect 117 135 120 137
rect 113 130 120 135
rect 113 128 115 130
rect 117 128 120 130
rect 113 126 120 128
rect 122 142 130 144
rect 122 140 125 142
rect 127 140 130 142
rect 122 133 130 140
rect 132 144 140 146
rect 132 142 135 144
rect 137 142 140 144
rect 132 137 140 142
rect 132 135 135 137
rect 137 135 140 137
rect 132 133 140 135
rect 142 144 149 146
rect 142 142 145 144
rect 147 142 149 144
rect 142 133 149 142
rect 122 126 128 133
rect 164 132 169 153
rect 162 130 169 132
rect 162 128 164 130
rect 166 128 169 130
rect 162 126 169 128
rect 171 151 183 153
rect 171 149 174 151
rect 176 149 183 151
rect 171 144 183 149
rect 200 144 205 153
rect 171 142 174 144
rect 176 142 185 144
rect 171 126 185 142
rect 187 137 195 144
rect 187 135 190 137
rect 192 135 195 137
rect 187 130 195 135
rect 187 128 190 130
rect 192 128 195 130
rect 187 126 195 128
rect 197 137 205 144
rect 197 135 200 137
rect 202 135 205 137
rect 197 126 205 135
rect 207 147 212 153
rect 207 145 214 147
rect 207 143 210 145
rect 212 143 214 145
rect 248 144 254 146
rect 207 141 214 143
rect 207 126 212 141
rect 239 139 244 144
rect 237 137 244 139
rect 237 135 239 137
rect 241 135 244 137
rect 237 130 244 135
rect 237 128 239 130
rect 241 128 244 130
rect 237 126 244 128
rect 246 142 254 144
rect 246 140 249 142
rect 251 140 254 142
rect 246 133 254 140
rect 256 144 264 146
rect 256 142 259 144
rect 261 142 264 144
rect 256 137 264 142
rect 256 135 259 137
rect 261 135 264 137
rect 256 133 264 135
rect 266 144 273 146
rect 266 142 269 144
rect 271 142 273 144
rect 266 133 273 142
rect 246 126 252 133
rect 288 132 293 153
rect 286 130 293 132
rect 286 128 288 130
rect 290 128 293 130
rect 286 126 293 128
rect 295 151 307 153
rect 295 149 298 151
rect 300 149 307 151
rect 295 144 307 149
rect 324 144 329 153
rect 295 142 298 144
rect 300 142 309 144
rect 295 126 309 142
rect 311 137 319 144
rect 311 135 314 137
rect 316 135 319 137
rect 311 130 319 135
rect 311 128 314 130
rect 316 128 319 130
rect 311 126 319 128
rect 321 137 329 144
rect 321 135 324 137
rect 326 135 329 137
rect 321 126 329 135
rect 331 147 336 153
rect 331 145 338 147
rect 331 143 334 145
rect 336 143 338 145
rect 331 141 338 143
rect 363 143 370 145
rect 363 141 365 143
rect 367 141 370 143
rect 331 126 336 141
rect 363 132 370 141
rect 372 143 380 145
rect 372 141 375 143
rect 377 141 380 143
rect 372 136 380 141
rect 372 134 375 136
rect 377 134 380 136
rect 372 132 380 134
rect 382 143 388 145
rect 403 143 410 145
rect 382 141 390 143
rect 382 139 385 141
rect 387 139 390 141
rect 382 132 390 139
rect 384 125 390 132
rect 392 138 397 143
rect 403 141 405 143
rect 407 141 410 143
rect 392 136 399 138
rect 392 134 395 136
rect 397 134 399 136
rect 392 129 399 134
rect 403 132 410 141
rect 412 143 420 145
rect 412 141 415 143
rect 417 141 420 143
rect 412 136 420 141
rect 412 134 415 136
rect 417 134 420 136
rect 412 132 420 134
rect 422 143 428 145
rect 452 146 457 152
rect 450 144 457 146
rect 422 141 430 143
rect 422 139 425 141
rect 427 139 430 141
rect 422 132 430 139
rect 392 127 395 129
rect 397 127 399 129
rect 392 125 399 127
rect 424 125 430 132
rect 432 138 437 143
rect 450 142 452 144
rect 454 142 457 144
rect 450 140 457 142
rect 432 136 439 138
rect 432 134 435 136
rect 437 134 439 136
rect 432 129 439 134
rect 432 127 435 129
rect 437 127 439 129
rect 432 125 439 127
rect 452 125 457 140
rect 459 143 464 152
rect 481 150 493 152
rect 481 148 488 150
rect 490 148 493 150
rect 481 143 493 148
rect 459 136 467 143
rect 459 134 462 136
rect 464 134 467 136
rect 459 125 467 134
rect 469 136 477 143
rect 469 134 472 136
rect 474 134 477 136
rect 469 129 477 134
rect 469 127 472 129
rect 474 127 477 129
rect 469 125 477 127
rect 479 141 488 143
rect 490 141 493 143
rect 479 125 493 141
rect 495 131 500 152
rect 515 143 522 145
rect 515 141 517 143
rect 519 141 522 143
rect 515 132 522 141
rect 524 143 532 145
rect 524 141 527 143
rect 529 141 532 143
rect 524 136 532 141
rect 524 134 527 136
rect 529 134 532 136
rect 524 132 532 134
rect 534 143 540 145
rect 568 143 575 145
rect 534 141 542 143
rect 534 139 537 141
rect 539 139 542 141
rect 534 132 542 139
rect 495 129 502 131
rect 495 127 498 129
rect 500 127 502 129
rect 495 125 502 127
rect 536 125 542 132
rect 544 138 549 143
rect 568 141 570 143
rect 572 141 575 143
rect 544 136 551 138
rect 544 134 547 136
rect 549 134 551 136
rect 544 129 551 134
rect 568 132 575 141
rect 577 143 585 145
rect 577 141 580 143
rect 582 141 585 143
rect 577 136 585 141
rect 577 134 580 136
rect 582 134 585 136
rect 577 132 585 134
rect 587 143 593 145
rect 608 143 615 145
rect 587 141 595 143
rect 587 139 590 141
rect 592 139 595 141
rect 587 132 595 139
rect 544 127 547 129
rect 549 127 551 129
rect 544 125 551 127
rect 589 125 595 132
rect 597 138 602 143
rect 608 141 610 143
rect 612 141 615 143
rect 597 136 604 138
rect 597 134 600 136
rect 602 134 604 136
rect 597 129 604 134
rect 608 132 615 141
rect 617 143 625 145
rect 617 141 620 143
rect 622 141 625 143
rect 617 136 625 141
rect 617 134 620 136
rect 622 134 625 136
rect 617 132 625 134
rect 627 143 633 145
rect 657 146 662 152
rect 655 144 662 146
rect 627 141 635 143
rect 627 139 630 141
rect 632 139 635 141
rect 627 132 635 139
rect 597 127 600 129
rect 602 127 604 129
rect 597 125 604 127
rect 629 125 635 132
rect 637 138 642 143
rect 655 142 657 144
rect 659 142 662 144
rect 655 140 662 142
rect 637 136 644 138
rect 637 134 640 136
rect 642 134 644 136
rect 637 129 644 134
rect 637 127 640 129
rect 642 127 644 129
rect 637 125 644 127
rect 657 125 662 140
rect 664 143 669 152
rect 686 150 698 152
rect 686 148 693 150
rect 695 148 698 150
rect 686 143 698 148
rect 664 136 672 143
rect 664 134 667 136
rect 669 134 672 136
rect 664 125 672 134
rect 674 136 682 143
rect 674 134 677 136
rect 679 134 682 136
rect 674 129 682 134
rect 674 127 677 129
rect 679 127 682 129
rect 674 125 682 127
rect 684 141 693 143
rect 695 141 698 143
rect 684 125 698 141
rect 700 131 705 152
rect 786 151 795 153
rect 786 149 788 151
rect 790 149 795 151
rect 720 143 727 145
rect 720 141 722 143
rect 724 141 727 143
rect 720 132 727 141
rect 729 143 737 145
rect 729 141 732 143
rect 734 141 737 143
rect 729 136 737 141
rect 729 134 732 136
rect 734 134 737 136
rect 729 132 737 134
rect 739 143 745 145
rect 786 143 795 149
rect 739 141 747 143
rect 739 139 742 141
rect 744 139 747 141
rect 739 132 747 139
rect 700 129 707 131
rect 700 127 703 129
rect 705 127 707 129
rect 700 125 707 127
rect 741 125 747 132
rect 749 138 754 143
rect 775 141 782 143
rect 775 139 777 141
rect 779 139 782 141
rect 749 136 756 138
rect 749 134 752 136
rect 754 134 756 136
rect 749 129 756 134
rect 775 134 782 139
rect 775 132 777 134
rect 779 132 782 134
rect 775 130 782 132
rect 749 127 752 129
rect 754 127 756 129
rect 749 125 756 127
rect 777 125 782 130
rect 784 132 795 143
rect 797 132 802 153
rect 804 146 809 153
rect 804 144 811 146
rect 826 144 832 146
rect 804 142 807 144
rect 809 142 811 144
rect 804 140 811 142
rect 804 132 809 140
rect 817 139 822 144
rect 815 137 822 139
rect 815 135 817 137
rect 819 135 822 137
rect 784 125 792 132
rect 815 130 822 135
rect 815 128 817 130
rect 819 128 822 130
rect 815 126 822 128
rect 824 142 832 144
rect 824 140 827 142
rect 829 140 832 142
rect 824 133 832 140
rect 834 144 842 146
rect 834 142 837 144
rect 839 142 842 144
rect 834 137 842 142
rect 834 135 837 137
rect 839 135 842 137
rect 834 133 842 135
rect 844 144 851 146
rect 844 142 847 144
rect 849 142 851 144
rect 844 133 851 142
rect 824 126 830 133
rect 866 132 871 153
rect 864 130 871 132
rect 864 128 866 130
rect 868 128 871 130
rect 864 126 871 128
rect 873 151 885 153
rect 873 149 876 151
rect 878 149 885 151
rect 873 144 885 149
rect 902 144 907 153
rect 873 142 876 144
rect 878 142 887 144
rect 873 126 887 142
rect 889 137 897 144
rect 889 135 892 137
rect 894 135 897 137
rect 889 130 897 135
rect 889 128 892 130
rect 894 128 897 130
rect 889 126 897 128
rect 899 137 907 144
rect 899 135 902 137
rect 904 135 907 137
rect 899 126 907 135
rect 909 147 914 153
rect 909 145 916 147
rect 909 143 912 145
rect 914 143 916 145
rect 931 144 937 146
rect 909 141 916 143
rect 909 126 914 141
rect 922 139 927 144
rect 920 137 927 139
rect 920 135 922 137
rect 924 135 927 137
rect 920 130 927 135
rect 920 128 922 130
rect 924 128 927 130
rect 920 126 927 128
rect 929 142 937 144
rect 929 140 932 142
rect 934 140 937 142
rect 929 133 937 140
rect 939 144 947 146
rect 939 142 942 144
rect 944 142 947 144
rect 939 137 947 142
rect 939 135 942 137
rect 944 135 947 137
rect 939 133 947 135
rect 949 144 956 146
rect 949 142 952 144
rect 954 142 956 144
rect 949 133 956 142
rect 929 126 935 133
rect 971 132 976 153
rect 969 130 976 132
rect 969 128 971 130
rect 973 128 976 130
rect 969 126 976 128
rect 978 151 990 153
rect 978 149 981 151
rect 983 149 990 151
rect 978 144 990 149
rect 1007 144 1012 153
rect 978 142 981 144
rect 983 142 992 144
rect 978 126 992 142
rect 994 137 1002 144
rect 994 135 997 137
rect 999 135 1002 137
rect 994 130 1002 135
rect 994 128 997 130
rect 999 128 1002 130
rect 994 126 1002 128
rect 1004 137 1012 144
rect 1004 135 1007 137
rect 1009 135 1012 137
rect 1004 126 1012 135
rect 1014 147 1019 153
rect 1036 151 1045 153
rect 1036 149 1038 151
rect 1040 149 1045 151
rect 1014 145 1021 147
rect 1014 143 1017 145
rect 1019 143 1021 145
rect 1036 143 1045 149
rect 1014 141 1021 143
rect 1025 141 1032 143
rect 1014 126 1019 141
rect 1025 139 1027 141
rect 1029 139 1032 141
rect 1025 134 1032 139
rect 1025 132 1027 134
rect 1029 132 1032 134
rect 1025 130 1032 132
rect 1027 125 1032 130
rect 1034 132 1045 143
rect 1047 132 1052 153
rect 1054 146 1059 153
rect 1054 144 1061 146
rect 1076 144 1082 146
rect 1054 142 1057 144
rect 1059 142 1061 144
rect 1054 140 1061 142
rect 1054 132 1059 140
rect 1067 139 1072 144
rect 1065 137 1072 139
rect 1065 135 1067 137
rect 1069 135 1072 137
rect 1034 125 1042 132
rect 1065 130 1072 135
rect 1065 128 1067 130
rect 1069 128 1072 130
rect 1065 126 1072 128
rect 1074 142 1082 144
rect 1074 140 1077 142
rect 1079 140 1082 142
rect 1074 133 1082 140
rect 1084 144 1092 146
rect 1084 142 1087 144
rect 1089 142 1092 144
rect 1084 137 1092 142
rect 1084 135 1087 137
rect 1089 135 1092 137
rect 1084 133 1092 135
rect 1094 144 1101 146
rect 1094 142 1097 144
rect 1099 142 1101 144
rect 1094 133 1101 142
rect 1074 126 1080 133
rect 1116 132 1121 153
rect 1114 130 1121 132
rect 1114 128 1116 130
rect 1118 128 1121 130
rect 1114 126 1121 128
rect 1123 151 1135 153
rect 1123 149 1126 151
rect 1128 149 1135 151
rect 1123 144 1135 149
rect 1152 144 1157 153
rect 1123 142 1126 144
rect 1128 142 1137 144
rect 1123 126 1137 142
rect 1139 137 1147 144
rect 1139 135 1142 137
rect 1144 135 1147 137
rect 1139 130 1147 135
rect 1139 128 1142 130
rect 1144 128 1147 130
rect 1139 126 1147 128
rect 1149 137 1157 144
rect 1149 135 1152 137
rect 1154 135 1157 137
rect 1149 126 1157 135
rect 1159 147 1164 153
rect 1159 145 1166 147
rect 1159 143 1162 145
rect 1164 143 1166 145
rect 1181 144 1187 146
rect 1159 141 1166 143
rect 1159 126 1164 141
rect 1172 139 1177 144
rect 1170 137 1177 139
rect 1170 135 1172 137
rect 1174 135 1177 137
rect 1170 130 1177 135
rect 1170 128 1172 130
rect 1174 128 1177 130
rect 1170 126 1177 128
rect 1179 142 1187 144
rect 1179 140 1182 142
rect 1184 140 1187 142
rect 1179 133 1187 140
rect 1189 144 1197 146
rect 1189 142 1192 144
rect 1194 142 1197 144
rect 1189 137 1197 142
rect 1189 135 1192 137
rect 1194 135 1197 137
rect 1189 133 1197 135
rect 1199 144 1206 146
rect 1199 142 1202 144
rect 1204 142 1206 144
rect 1199 133 1206 142
rect 1179 126 1185 133
rect 1221 132 1226 153
rect 1219 130 1226 132
rect 1219 128 1221 130
rect 1223 128 1226 130
rect 1219 126 1226 128
rect 1228 151 1240 153
rect 1228 149 1231 151
rect 1233 149 1240 151
rect 1228 144 1240 149
rect 1257 144 1262 153
rect 1228 142 1231 144
rect 1233 142 1242 144
rect 1228 126 1242 142
rect 1244 137 1252 144
rect 1244 135 1247 137
rect 1249 135 1252 137
rect 1244 130 1252 135
rect 1244 128 1247 130
rect 1249 128 1252 130
rect 1244 126 1252 128
rect 1254 137 1262 144
rect 1254 135 1257 137
rect 1259 135 1262 137
rect 1254 126 1262 135
rect 1264 147 1269 153
rect 1286 151 1295 153
rect 1286 149 1288 151
rect 1290 149 1295 151
rect 1264 145 1271 147
rect 1264 143 1267 145
rect 1269 143 1271 145
rect 1286 143 1295 149
rect 1264 141 1271 143
rect 1275 141 1282 143
rect 1264 126 1269 141
rect 1275 139 1277 141
rect 1279 139 1282 141
rect 1275 134 1282 139
rect 1275 132 1277 134
rect 1279 132 1282 134
rect 1275 130 1282 132
rect 1277 125 1282 130
rect 1284 132 1295 143
rect 1297 132 1302 153
rect 1304 146 1309 153
rect 1304 144 1311 146
rect 1326 144 1332 146
rect 1304 142 1307 144
rect 1309 142 1311 144
rect 1304 140 1311 142
rect 1304 132 1309 140
rect 1317 139 1322 144
rect 1315 137 1322 139
rect 1315 135 1317 137
rect 1319 135 1322 137
rect 1284 125 1292 132
rect 1315 130 1322 135
rect 1315 128 1317 130
rect 1319 128 1322 130
rect 1315 126 1322 128
rect 1324 142 1332 144
rect 1324 140 1327 142
rect 1329 140 1332 142
rect 1324 133 1332 140
rect 1334 144 1342 146
rect 1334 142 1337 144
rect 1339 142 1342 144
rect 1334 137 1342 142
rect 1334 135 1337 137
rect 1339 135 1342 137
rect 1334 133 1342 135
rect 1344 144 1351 146
rect 1344 142 1347 144
rect 1349 142 1351 144
rect 1344 133 1351 142
rect 1324 126 1330 133
rect 1366 132 1371 153
rect 1364 130 1371 132
rect 1364 128 1366 130
rect 1368 128 1371 130
rect 1364 126 1371 128
rect 1373 151 1385 153
rect 1373 149 1376 151
rect 1378 149 1385 151
rect 1373 144 1385 149
rect 1402 144 1407 153
rect 1373 142 1376 144
rect 1378 142 1387 144
rect 1373 126 1387 142
rect 1389 137 1397 144
rect 1389 135 1392 137
rect 1394 135 1397 137
rect 1389 130 1397 135
rect 1389 128 1392 130
rect 1394 128 1397 130
rect 1389 126 1397 128
rect 1399 137 1407 144
rect 1399 135 1402 137
rect 1404 135 1407 137
rect 1399 126 1407 135
rect 1409 147 1414 153
rect 1409 145 1416 147
rect 1409 143 1412 145
rect 1414 143 1416 145
rect 1431 144 1437 146
rect 1409 141 1416 143
rect 1409 126 1414 141
rect 1422 139 1427 144
rect 1420 137 1427 139
rect 1420 135 1422 137
rect 1424 135 1427 137
rect 1420 130 1427 135
rect 1420 128 1422 130
rect 1424 128 1427 130
rect 1420 126 1427 128
rect 1429 142 1437 144
rect 1429 140 1432 142
rect 1434 140 1437 142
rect 1429 133 1437 140
rect 1439 144 1447 146
rect 1439 142 1442 144
rect 1444 142 1447 144
rect 1439 137 1447 142
rect 1439 135 1442 137
rect 1444 135 1447 137
rect 1439 133 1447 135
rect 1449 144 1456 146
rect 1449 142 1452 144
rect 1454 142 1456 144
rect 1449 133 1456 142
rect 1429 126 1435 133
rect 1471 132 1476 153
rect 1469 130 1476 132
rect 1469 128 1471 130
rect 1473 128 1476 130
rect 1469 126 1476 128
rect 1478 151 1490 153
rect 1478 149 1481 151
rect 1483 149 1490 151
rect 1478 144 1490 149
rect 1507 144 1512 153
rect 1478 142 1481 144
rect 1483 142 1492 144
rect 1478 126 1492 142
rect 1494 137 1502 144
rect 1494 135 1497 137
rect 1499 135 1502 137
rect 1494 130 1502 135
rect 1494 128 1497 130
rect 1499 128 1502 130
rect 1494 126 1502 128
rect 1504 137 1512 144
rect 1504 135 1507 137
rect 1509 135 1512 137
rect 1504 126 1512 135
rect 1514 147 1519 153
rect 1536 151 1545 153
rect 1536 149 1538 151
rect 1540 149 1545 151
rect 1514 145 1521 147
rect 1514 143 1517 145
rect 1519 143 1521 145
rect 1536 143 1545 149
rect 1514 141 1521 143
rect 1525 141 1532 143
rect 1514 126 1519 141
rect 1525 139 1527 141
rect 1529 139 1532 141
rect 1525 134 1532 139
rect 1525 132 1527 134
rect 1529 132 1532 134
rect 1525 130 1532 132
rect 1527 125 1532 130
rect 1534 132 1545 143
rect 1547 132 1552 153
rect 1554 146 1559 153
rect 1554 144 1561 146
rect 1576 144 1582 146
rect 1554 142 1557 144
rect 1559 142 1561 144
rect 1554 140 1561 142
rect 1554 132 1559 140
rect 1567 139 1572 144
rect 1565 137 1572 139
rect 1565 135 1567 137
rect 1569 135 1572 137
rect 1534 125 1542 132
rect 1565 130 1572 135
rect 1565 128 1567 130
rect 1569 128 1572 130
rect 1565 126 1572 128
rect 1574 142 1582 144
rect 1574 140 1577 142
rect 1579 140 1582 142
rect 1574 133 1582 140
rect 1584 144 1592 146
rect 1584 142 1587 144
rect 1589 142 1592 144
rect 1584 137 1592 142
rect 1584 135 1587 137
rect 1589 135 1592 137
rect 1584 133 1592 135
rect 1594 144 1601 146
rect 1594 142 1597 144
rect 1599 142 1601 144
rect 1594 133 1601 142
rect 1574 126 1580 133
rect 1616 132 1621 153
rect 1614 130 1621 132
rect 1614 128 1616 130
rect 1618 128 1621 130
rect 1614 126 1621 128
rect 1623 151 1635 153
rect 1623 149 1626 151
rect 1628 149 1635 151
rect 1623 144 1635 149
rect 1652 144 1657 153
rect 1623 142 1626 144
rect 1628 142 1637 144
rect 1623 126 1637 142
rect 1639 137 1647 144
rect 1639 135 1642 137
rect 1644 135 1647 137
rect 1639 130 1647 135
rect 1639 128 1642 130
rect 1644 128 1647 130
rect 1639 126 1647 128
rect 1649 137 1657 144
rect 1649 135 1652 137
rect 1654 135 1657 137
rect 1649 126 1657 135
rect 1659 147 1664 153
rect 1659 145 1666 147
rect 1659 143 1662 145
rect 1664 143 1666 145
rect 1681 144 1687 146
rect 1659 141 1666 143
rect 1659 126 1664 141
rect 1672 139 1677 144
rect 1670 137 1677 139
rect 1670 135 1672 137
rect 1674 135 1677 137
rect 1670 130 1677 135
rect 1670 128 1672 130
rect 1674 128 1677 130
rect 1670 126 1677 128
rect 1679 142 1687 144
rect 1679 140 1682 142
rect 1684 140 1687 142
rect 1679 133 1687 140
rect 1689 144 1697 146
rect 1689 142 1692 144
rect 1694 142 1697 144
rect 1689 137 1697 142
rect 1689 135 1692 137
rect 1694 135 1697 137
rect 1689 133 1697 135
rect 1699 144 1706 146
rect 1699 142 1702 144
rect 1704 142 1706 144
rect 1699 133 1706 142
rect 1679 126 1685 133
rect 1721 132 1726 153
rect 1719 130 1726 132
rect 1719 128 1721 130
rect 1723 128 1726 130
rect 1719 126 1726 128
rect 1728 151 1740 153
rect 1728 149 1731 151
rect 1733 149 1740 151
rect 1728 144 1740 149
rect 1757 144 1762 153
rect 1728 142 1731 144
rect 1733 142 1742 144
rect 1728 126 1742 142
rect 1744 137 1752 144
rect 1744 135 1747 137
rect 1749 135 1752 137
rect 1744 130 1752 135
rect 1744 128 1747 130
rect 1749 128 1752 130
rect 1744 126 1752 128
rect 1754 137 1762 144
rect 1754 135 1757 137
rect 1759 135 1762 137
rect 1754 126 1762 135
rect 1764 147 1769 153
rect 1764 145 1771 147
rect 1764 143 1767 145
rect 1769 143 1771 145
rect 1834 144 1840 146
rect 1764 141 1771 143
rect 1764 126 1769 141
rect 1825 139 1830 144
rect 1823 137 1830 139
rect 1823 135 1825 137
rect 1827 135 1830 137
rect 1823 130 1830 135
rect 1823 128 1825 130
rect 1827 128 1830 130
rect 1823 126 1830 128
rect 1832 142 1840 144
rect 1832 140 1835 142
rect 1837 140 1840 142
rect 1832 133 1840 140
rect 1842 144 1850 146
rect 1842 142 1845 144
rect 1847 142 1850 144
rect 1842 137 1850 142
rect 1842 135 1845 137
rect 1847 135 1850 137
rect 1842 133 1850 135
rect 1852 144 1859 146
rect 1852 142 1855 144
rect 1857 142 1859 144
rect 1852 133 1859 142
rect 1863 144 1870 146
rect 1863 142 1865 144
rect 1867 142 1870 144
rect 1863 133 1870 142
rect 1872 144 1880 146
rect 1872 142 1875 144
rect 1877 142 1880 144
rect 1872 137 1880 142
rect 1872 135 1875 137
rect 1877 135 1880 137
rect 1872 133 1880 135
rect 1882 144 1888 146
rect 1914 144 1920 146
rect 1882 142 1890 144
rect 1882 140 1885 142
rect 1887 140 1890 142
rect 1882 133 1890 140
rect 1832 126 1838 133
rect 1884 126 1890 133
rect 1892 139 1897 144
rect 1905 139 1910 144
rect 1892 137 1899 139
rect 1892 135 1895 137
rect 1897 135 1899 137
rect 1892 130 1899 135
rect 1892 128 1895 130
rect 1897 128 1899 130
rect 1892 126 1899 128
rect 1903 137 1910 139
rect 1903 135 1905 137
rect 1907 135 1910 137
rect 1903 130 1910 135
rect 1903 128 1905 130
rect 1907 128 1910 130
rect 1903 126 1910 128
rect 1912 142 1920 144
rect 1912 140 1915 142
rect 1917 140 1920 142
rect 1912 133 1920 140
rect 1922 144 1930 146
rect 1922 142 1925 144
rect 1927 142 1930 144
rect 1922 137 1930 142
rect 1922 135 1925 137
rect 1927 135 1930 137
rect 1922 133 1930 135
rect 1932 144 1939 146
rect 1932 142 1935 144
rect 1937 142 1939 144
rect 1932 133 1939 142
rect 1912 126 1918 133
rect 1954 132 1959 153
rect 1952 130 1959 132
rect 1952 128 1954 130
rect 1956 128 1959 130
rect 1952 126 1959 128
rect 1961 151 1973 153
rect 1961 149 1964 151
rect 1966 149 1973 151
rect 1961 144 1973 149
rect 1990 144 1995 153
rect 1961 142 1964 144
rect 1966 142 1975 144
rect 1961 126 1975 142
rect 1977 137 1985 144
rect 1977 135 1980 137
rect 1982 135 1985 137
rect 1977 130 1985 135
rect 1977 128 1980 130
rect 1982 128 1985 130
rect 1977 126 1985 128
rect 1987 137 1995 144
rect 1987 135 1990 137
rect 1992 135 1995 137
rect 1987 126 1995 135
rect 1997 147 2002 153
rect 1997 145 2004 147
rect 1997 143 2000 145
rect 2002 143 2004 145
rect 1997 141 2004 143
rect 1997 126 2002 141
rect 9 34 14 39
rect 7 32 14 34
rect 7 30 9 32
rect 11 30 14 32
rect 7 25 14 30
rect 7 23 9 25
rect 11 23 14 25
rect 7 21 14 23
rect 16 32 24 39
rect 47 36 54 38
rect 47 34 49 36
rect 51 34 54 36
rect 16 21 27 32
rect 18 15 27 21
rect 18 13 20 15
rect 22 13 27 15
rect 18 11 27 13
rect 29 11 34 32
rect 36 24 41 32
rect 47 29 54 34
rect 47 27 49 29
rect 51 27 54 29
rect 47 25 54 27
rect 36 22 43 24
rect 36 20 39 22
rect 41 20 43 22
rect 49 20 54 25
rect 56 31 62 38
rect 96 36 103 38
rect 96 34 98 36
rect 100 34 103 36
rect 96 32 103 34
rect 56 24 64 31
rect 56 22 59 24
rect 61 22 64 24
rect 56 20 64 22
rect 36 18 43 20
rect 36 11 41 18
rect 58 18 64 20
rect 66 29 74 31
rect 66 27 69 29
rect 71 27 74 29
rect 66 22 74 27
rect 66 20 69 22
rect 71 20 74 22
rect 66 18 74 20
rect 76 22 83 31
rect 76 20 79 22
rect 81 20 83 22
rect 76 18 83 20
rect 98 11 103 32
rect 105 22 119 38
rect 105 20 108 22
rect 110 20 119 22
rect 121 36 129 38
rect 121 34 124 36
rect 126 34 129 36
rect 121 29 129 34
rect 121 27 124 29
rect 126 27 129 29
rect 121 20 129 27
rect 131 29 139 38
rect 131 27 134 29
rect 136 27 139 29
rect 131 20 139 27
rect 105 15 117 20
rect 105 13 108 15
rect 110 13 117 15
rect 105 11 117 13
rect 134 11 139 20
rect 141 23 146 38
rect 152 36 159 38
rect 152 34 154 36
rect 156 34 159 36
rect 152 29 159 34
rect 152 27 154 29
rect 156 27 159 29
rect 152 25 159 27
rect 141 21 148 23
rect 141 19 144 21
rect 146 19 148 21
rect 154 20 159 25
rect 161 31 167 38
rect 201 36 208 38
rect 201 34 203 36
rect 205 34 208 36
rect 201 32 208 34
rect 161 24 169 31
rect 161 22 164 24
rect 166 22 169 24
rect 161 20 169 22
rect 141 17 148 19
rect 141 11 146 17
rect 163 18 169 20
rect 171 29 179 31
rect 171 27 174 29
rect 176 27 179 29
rect 171 22 179 27
rect 171 20 174 22
rect 176 20 179 22
rect 171 18 179 20
rect 181 22 188 31
rect 181 20 184 22
rect 186 20 188 22
rect 181 18 188 20
rect 203 11 208 32
rect 210 22 224 38
rect 210 20 213 22
rect 215 20 224 22
rect 226 36 234 38
rect 226 34 229 36
rect 231 34 234 36
rect 226 29 234 34
rect 226 27 229 29
rect 231 27 234 29
rect 226 20 234 27
rect 236 29 244 38
rect 236 27 239 29
rect 241 27 244 29
rect 236 20 244 27
rect 210 15 222 20
rect 210 13 213 15
rect 215 13 222 15
rect 210 11 222 13
rect 239 11 244 20
rect 246 23 251 38
rect 259 34 264 39
rect 257 32 264 34
rect 257 30 259 32
rect 261 30 264 32
rect 257 25 264 30
rect 257 23 259 25
rect 261 23 264 25
rect 246 21 253 23
rect 257 21 264 23
rect 266 32 274 39
rect 297 36 304 38
rect 297 34 299 36
rect 301 34 304 36
rect 266 21 277 32
rect 246 19 249 21
rect 251 19 253 21
rect 246 17 253 19
rect 246 11 251 17
rect 268 15 277 21
rect 268 13 270 15
rect 272 13 277 15
rect 268 11 277 13
rect 279 11 284 32
rect 286 24 291 32
rect 297 29 304 34
rect 297 27 299 29
rect 301 27 304 29
rect 297 25 304 27
rect 286 22 293 24
rect 286 20 289 22
rect 291 20 293 22
rect 299 20 304 25
rect 306 31 312 38
rect 346 36 353 38
rect 346 34 348 36
rect 350 34 353 36
rect 346 32 353 34
rect 306 24 314 31
rect 306 22 309 24
rect 311 22 314 24
rect 306 20 314 22
rect 286 18 293 20
rect 286 11 291 18
rect 308 18 314 20
rect 316 29 324 31
rect 316 27 319 29
rect 321 27 324 29
rect 316 22 324 27
rect 316 20 319 22
rect 321 20 324 22
rect 316 18 324 20
rect 326 22 333 31
rect 326 20 329 22
rect 331 20 333 22
rect 326 18 333 20
rect 348 11 353 32
rect 355 22 369 38
rect 355 20 358 22
rect 360 20 369 22
rect 371 36 379 38
rect 371 34 374 36
rect 376 34 379 36
rect 371 29 379 34
rect 371 27 374 29
rect 376 27 379 29
rect 371 20 379 27
rect 381 29 389 38
rect 381 27 384 29
rect 386 27 389 29
rect 381 20 389 27
rect 355 15 367 20
rect 355 13 358 15
rect 360 13 367 15
rect 355 11 367 13
rect 384 11 389 20
rect 391 23 396 38
rect 402 36 409 38
rect 402 34 404 36
rect 406 34 409 36
rect 402 29 409 34
rect 402 27 404 29
rect 406 27 409 29
rect 402 25 409 27
rect 391 21 398 23
rect 391 19 394 21
rect 396 19 398 21
rect 404 20 409 25
rect 411 31 417 38
rect 451 36 458 38
rect 451 34 453 36
rect 455 34 458 36
rect 451 32 458 34
rect 411 24 419 31
rect 411 22 414 24
rect 416 22 419 24
rect 411 20 419 22
rect 391 17 398 19
rect 391 11 396 17
rect 413 18 419 20
rect 421 29 429 31
rect 421 27 424 29
rect 426 27 429 29
rect 421 22 429 27
rect 421 20 424 22
rect 426 20 429 22
rect 421 18 429 20
rect 431 22 438 31
rect 431 20 434 22
rect 436 20 438 22
rect 431 18 438 20
rect 453 11 458 32
rect 460 22 474 38
rect 460 20 463 22
rect 465 20 474 22
rect 476 36 484 38
rect 476 34 479 36
rect 481 34 484 36
rect 476 29 484 34
rect 476 27 479 29
rect 481 27 484 29
rect 476 20 484 27
rect 486 29 494 38
rect 486 27 489 29
rect 491 27 494 29
rect 486 20 494 27
rect 460 15 472 20
rect 460 13 463 15
rect 465 13 472 15
rect 460 11 472 13
rect 489 11 494 20
rect 496 23 501 38
rect 509 34 514 39
rect 507 32 514 34
rect 507 30 509 32
rect 511 30 514 32
rect 507 25 514 30
rect 507 23 509 25
rect 511 23 514 25
rect 496 21 503 23
rect 507 21 514 23
rect 516 32 524 39
rect 547 36 554 38
rect 547 34 549 36
rect 551 34 554 36
rect 516 21 527 32
rect 496 19 499 21
rect 501 19 503 21
rect 496 17 503 19
rect 496 11 501 17
rect 518 15 527 21
rect 518 13 520 15
rect 522 13 527 15
rect 518 11 527 13
rect 529 11 534 32
rect 536 24 541 32
rect 547 29 554 34
rect 547 27 549 29
rect 551 27 554 29
rect 547 25 554 27
rect 536 22 543 24
rect 536 20 539 22
rect 541 20 543 22
rect 549 20 554 25
rect 556 31 562 38
rect 596 36 603 38
rect 596 34 598 36
rect 600 34 603 36
rect 596 32 603 34
rect 556 24 564 31
rect 556 22 559 24
rect 561 22 564 24
rect 556 20 564 22
rect 536 18 543 20
rect 536 11 541 18
rect 558 18 564 20
rect 566 29 574 31
rect 566 27 569 29
rect 571 27 574 29
rect 566 22 574 27
rect 566 20 569 22
rect 571 20 574 22
rect 566 18 574 20
rect 576 22 583 31
rect 576 20 579 22
rect 581 20 583 22
rect 576 18 583 20
rect 598 11 603 32
rect 605 22 619 38
rect 605 20 608 22
rect 610 20 619 22
rect 621 36 629 38
rect 621 34 624 36
rect 626 34 629 36
rect 621 29 629 34
rect 621 27 624 29
rect 626 27 629 29
rect 621 20 629 27
rect 631 29 639 38
rect 631 27 634 29
rect 636 27 639 29
rect 631 20 639 27
rect 605 15 617 20
rect 605 13 608 15
rect 610 13 617 15
rect 605 11 617 13
rect 634 11 639 20
rect 641 23 646 38
rect 652 36 659 38
rect 652 34 654 36
rect 656 34 659 36
rect 652 29 659 34
rect 652 27 654 29
rect 656 27 659 29
rect 652 25 659 27
rect 641 21 648 23
rect 641 19 644 21
rect 646 19 648 21
rect 654 20 659 25
rect 661 31 667 38
rect 701 36 708 38
rect 701 34 703 36
rect 705 34 708 36
rect 701 32 708 34
rect 661 24 669 31
rect 661 22 664 24
rect 666 22 669 24
rect 661 20 669 22
rect 641 17 648 19
rect 641 11 646 17
rect 663 18 669 20
rect 671 29 679 31
rect 671 27 674 29
rect 676 27 679 29
rect 671 22 679 27
rect 671 20 674 22
rect 676 20 679 22
rect 671 18 679 20
rect 681 22 688 31
rect 681 20 684 22
rect 686 20 688 22
rect 681 18 688 20
rect 703 11 708 32
rect 710 22 724 38
rect 710 20 713 22
rect 715 20 724 22
rect 726 36 734 38
rect 726 34 729 36
rect 731 34 734 36
rect 726 29 734 34
rect 726 27 729 29
rect 731 27 734 29
rect 726 20 734 27
rect 736 29 744 38
rect 736 27 739 29
rect 741 27 744 29
rect 736 20 744 27
rect 710 15 722 20
rect 710 13 713 15
rect 715 13 722 15
rect 710 11 722 13
rect 739 11 744 20
rect 746 23 751 38
rect 759 34 764 39
rect 757 32 764 34
rect 757 30 759 32
rect 761 30 764 32
rect 757 25 764 30
rect 757 23 759 25
rect 761 23 764 25
rect 746 21 753 23
rect 757 21 764 23
rect 766 32 774 39
rect 797 36 804 38
rect 797 34 799 36
rect 801 34 804 36
rect 766 21 777 32
rect 746 19 749 21
rect 751 19 753 21
rect 746 17 753 19
rect 746 11 751 17
rect 768 15 777 21
rect 768 13 770 15
rect 772 13 777 15
rect 768 11 777 13
rect 779 11 784 32
rect 786 24 791 32
rect 797 29 804 34
rect 797 27 799 29
rect 801 27 804 29
rect 797 25 804 27
rect 786 22 793 24
rect 786 20 789 22
rect 791 20 793 22
rect 799 20 804 25
rect 806 31 812 38
rect 846 36 853 38
rect 846 34 848 36
rect 850 34 853 36
rect 846 32 853 34
rect 806 24 814 31
rect 806 22 809 24
rect 811 22 814 24
rect 806 20 814 22
rect 786 18 793 20
rect 786 11 791 18
rect 808 18 814 20
rect 816 29 824 31
rect 816 27 819 29
rect 821 27 824 29
rect 816 22 824 27
rect 816 20 819 22
rect 821 20 824 22
rect 816 18 824 20
rect 826 22 833 31
rect 826 20 829 22
rect 831 20 833 22
rect 826 18 833 20
rect 848 11 853 32
rect 855 22 869 38
rect 855 20 858 22
rect 860 20 869 22
rect 871 36 879 38
rect 871 34 874 36
rect 876 34 879 36
rect 871 29 879 34
rect 871 27 874 29
rect 876 27 879 29
rect 871 20 879 27
rect 881 29 889 38
rect 881 27 884 29
rect 886 27 889 29
rect 881 20 889 27
rect 855 15 867 20
rect 855 13 858 15
rect 860 13 867 15
rect 855 11 867 13
rect 884 11 889 20
rect 891 23 896 38
rect 902 36 909 38
rect 902 34 904 36
rect 906 34 909 36
rect 902 29 909 34
rect 902 27 904 29
rect 906 27 909 29
rect 902 25 909 27
rect 891 21 898 23
rect 891 19 894 21
rect 896 19 898 21
rect 904 20 909 25
rect 911 31 917 38
rect 951 36 958 38
rect 951 34 953 36
rect 955 34 958 36
rect 951 32 958 34
rect 911 24 919 31
rect 911 22 914 24
rect 916 22 919 24
rect 911 20 919 22
rect 891 17 898 19
rect 891 11 896 17
rect 913 18 919 20
rect 921 29 929 31
rect 921 27 924 29
rect 926 27 929 29
rect 921 22 929 27
rect 921 20 924 22
rect 926 20 929 22
rect 921 18 929 20
rect 931 22 938 31
rect 931 20 934 22
rect 936 20 938 22
rect 931 18 938 20
rect 953 11 958 32
rect 960 22 974 38
rect 960 20 963 22
rect 965 20 974 22
rect 976 36 984 38
rect 976 34 979 36
rect 981 34 984 36
rect 976 29 984 34
rect 976 27 979 29
rect 981 27 984 29
rect 976 20 984 27
rect 986 29 994 38
rect 986 27 989 29
rect 991 27 994 29
rect 986 20 994 27
rect 960 15 972 20
rect 960 13 963 15
rect 965 13 972 15
rect 960 11 972 13
rect 989 11 994 20
rect 996 23 1001 38
rect 1019 34 1024 39
rect 1017 32 1024 34
rect 1017 30 1019 32
rect 1021 30 1024 32
rect 1017 25 1024 30
rect 1017 23 1019 25
rect 1021 23 1024 25
rect 996 21 1003 23
rect 1017 21 1024 23
rect 1026 32 1034 39
rect 1057 36 1064 38
rect 1057 34 1059 36
rect 1061 34 1064 36
rect 1026 21 1037 32
rect 996 19 999 21
rect 1001 19 1003 21
rect 996 17 1003 19
rect 996 11 1001 17
rect 1028 15 1037 21
rect 1028 13 1030 15
rect 1032 13 1037 15
rect 1028 11 1037 13
rect 1039 11 1044 32
rect 1046 24 1051 32
rect 1057 29 1064 34
rect 1057 27 1059 29
rect 1061 27 1064 29
rect 1057 25 1064 27
rect 1046 22 1053 24
rect 1046 20 1049 22
rect 1051 20 1053 22
rect 1059 20 1064 25
rect 1066 31 1072 38
rect 1106 36 1113 38
rect 1106 34 1108 36
rect 1110 34 1113 36
rect 1106 32 1113 34
rect 1066 24 1074 31
rect 1066 22 1069 24
rect 1071 22 1074 24
rect 1066 20 1074 22
rect 1046 18 1053 20
rect 1046 11 1051 18
rect 1068 18 1074 20
rect 1076 29 1084 31
rect 1076 27 1079 29
rect 1081 27 1084 29
rect 1076 22 1084 27
rect 1076 20 1079 22
rect 1081 20 1084 22
rect 1076 18 1084 20
rect 1086 22 1093 31
rect 1086 20 1089 22
rect 1091 20 1093 22
rect 1086 18 1093 20
rect 1108 11 1113 32
rect 1115 22 1129 38
rect 1115 20 1118 22
rect 1120 20 1129 22
rect 1131 36 1139 38
rect 1131 34 1134 36
rect 1136 34 1139 36
rect 1131 29 1139 34
rect 1131 27 1134 29
rect 1136 27 1139 29
rect 1131 20 1139 27
rect 1141 29 1149 38
rect 1141 27 1144 29
rect 1146 27 1149 29
rect 1141 20 1149 27
rect 1115 15 1127 20
rect 1115 13 1118 15
rect 1120 13 1127 15
rect 1115 11 1127 13
rect 1144 11 1149 20
rect 1151 23 1156 38
rect 1162 36 1169 38
rect 1162 34 1164 36
rect 1166 34 1169 36
rect 1162 29 1169 34
rect 1162 27 1164 29
rect 1166 27 1169 29
rect 1162 25 1169 27
rect 1151 21 1158 23
rect 1151 19 1154 21
rect 1156 19 1158 21
rect 1164 20 1169 25
rect 1171 31 1177 38
rect 1211 36 1218 38
rect 1211 34 1213 36
rect 1215 34 1218 36
rect 1211 32 1218 34
rect 1171 24 1179 31
rect 1171 22 1174 24
rect 1176 22 1179 24
rect 1171 20 1179 22
rect 1151 17 1158 19
rect 1151 11 1156 17
rect 1173 18 1179 20
rect 1181 29 1189 31
rect 1181 27 1184 29
rect 1186 27 1189 29
rect 1181 22 1189 27
rect 1181 20 1184 22
rect 1186 20 1189 22
rect 1181 18 1189 20
rect 1191 22 1198 31
rect 1191 20 1194 22
rect 1196 20 1198 22
rect 1191 18 1198 20
rect 1213 11 1218 32
rect 1220 22 1234 38
rect 1220 20 1223 22
rect 1225 20 1234 22
rect 1236 36 1244 38
rect 1236 34 1239 36
rect 1241 34 1244 36
rect 1236 29 1244 34
rect 1236 27 1239 29
rect 1241 27 1244 29
rect 1236 20 1244 27
rect 1246 29 1254 38
rect 1246 27 1249 29
rect 1251 27 1254 29
rect 1246 20 1254 27
rect 1220 15 1232 20
rect 1220 13 1223 15
rect 1225 13 1232 15
rect 1220 11 1232 13
rect 1249 11 1254 20
rect 1256 23 1261 38
rect 1269 34 1274 39
rect 1267 32 1274 34
rect 1267 30 1269 32
rect 1271 30 1274 32
rect 1267 25 1274 30
rect 1267 23 1269 25
rect 1271 23 1274 25
rect 1256 21 1263 23
rect 1267 21 1274 23
rect 1276 32 1284 39
rect 1307 36 1314 38
rect 1307 34 1309 36
rect 1311 34 1314 36
rect 1276 21 1287 32
rect 1256 19 1259 21
rect 1261 19 1263 21
rect 1256 17 1263 19
rect 1256 11 1261 17
rect 1278 15 1287 21
rect 1278 13 1280 15
rect 1282 13 1287 15
rect 1278 11 1287 13
rect 1289 11 1294 32
rect 1296 24 1301 32
rect 1307 29 1314 34
rect 1307 27 1309 29
rect 1311 27 1314 29
rect 1307 25 1314 27
rect 1296 22 1303 24
rect 1296 20 1299 22
rect 1301 20 1303 22
rect 1309 20 1314 25
rect 1316 31 1322 38
rect 1356 36 1363 38
rect 1356 34 1358 36
rect 1360 34 1363 36
rect 1356 32 1363 34
rect 1316 24 1324 31
rect 1316 22 1319 24
rect 1321 22 1324 24
rect 1316 20 1324 22
rect 1296 18 1303 20
rect 1296 11 1301 18
rect 1318 18 1324 20
rect 1326 29 1334 31
rect 1326 27 1329 29
rect 1331 27 1334 29
rect 1326 22 1334 27
rect 1326 20 1329 22
rect 1331 20 1334 22
rect 1326 18 1334 20
rect 1336 22 1343 31
rect 1336 20 1339 22
rect 1341 20 1343 22
rect 1336 18 1343 20
rect 1358 11 1363 32
rect 1365 22 1379 38
rect 1365 20 1368 22
rect 1370 20 1379 22
rect 1381 36 1389 38
rect 1381 34 1384 36
rect 1386 34 1389 36
rect 1381 29 1389 34
rect 1381 27 1384 29
rect 1386 27 1389 29
rect 1381 20 1389 27
rect 1391 29 1399 38
rect 1391 27 1394 29
rect 1396 27 1399 29
rect 1391 20 1399 27
rect 1365 15 1377 20
rect 1365 13 1368 15
rect 1370 13 1377 15
rect 1365 11 1377 13
rect 1394 11 1399 20
rect 1401 23 1406 38
rect 1412 36 1419 38
rect 1412 34 1414 36
rect 1416 34 1419 36
rect 1412 29 1419 34
rect 1412 27 1414 29
rect 1416 27 1419 29
rect 1412 25 1419 27
rect 1401 21 1408 23
rect 1401 19 1404 21
rect 1406 19 1408 21
rect 1414 20 1419 25
rect 1421 31 1427 38
rect 1461 36 1468 38
rect 1461 34 1463 36
rect 1465 34 1468 36
rect 1461 32 1468 34
rect 1421 24 1429 31
rect 1421 22 1424 24
rect 1426 22 1429 24
rect 1421 20 1429 22
rect 1401 17 1408 19
rect 1401 11 1406 17
rect 1423 18 1429 20
rect 1431 29 1439 31
rect 1431 27 1434 29
rect 1436 27 1439 29
rect 1431 22 1439 27
rect 1431 20 1434 22
rect 1436 20 1439 22
rect 1431 18 1439 20
rect 1441 22 1448 31
rect 1441 20 1444 22
rect 1446 20 1448 22
rect 1441 18 1448 20
rect 1463 11 1468 32
rect 1470 22 1484 38
rect 1470 20 1473 22
rect 1475 20 1484 22
rect 1486 36 1494 38
rect 1486 34 1489 36
rect 1491 34 1494 36
rect 1486 29 1494 34
rect 1486 27 1489 29
rect 1491 27 1494 29
rect 1486 20 1494 27
rect 1496 29 1504 38
rect 1496 27 1499 29
rect 1501 27 1504 29
rect 1496 20 1504 27
rect 1470 15 1482 20
rect 1470 13 1473 15
rect 1475 13 1482 15
rect 1470 11 1482 13
rect 1499 11 1504 20
rect 1506 23 1511 38
rect 1519 34 1524 39
rect 1517 32 1524 34
rect 1517 30 1519 32
rect 1521 30 1524 32
rect 1517 25 1524 30
rect 1517 23 1519 25
rect 1521 23 1524 25
rect 1506 21 1513 23
rect 1517 21 1524 23
rect 1526 32 1534 39
rect 1557 36 1564 38
rect 1557 34 1559 36
rect 1561 34 1564 36
rect 1526 21 1537 32
rect 1506 19 1509 21
rect 1511 19 1513 21
rect 1506 17 1513 19
rect 1506 11 1511 17
rect 1528 15 1537 21
rect 1528 13 1530 15
rect 1532 13 1537 15
rect 1528 11 1537 13
rect 1539 11 1544 32
rect 1546 24 1551 32
rect 1557 29 1564 34
rect 1557 27 1559 29
rect 1561 27 1564 29
rect 1557 25 1564 27
rect 1546 22 1553 24
rect 1546 20 1549 22
rect 1551 20 1553 22
rect 1559 20 1564 25
rect 1566 31 1572 38
rect 1606 36 1613 38
rect 1606 34 1608 36
rect 1610 34 1613 36
rect 1606 32 1613 34
rect 1566 24 1574 31
rect 1566 22 1569 24
rect 1571 22 1574 24
rect 1566 20 1574 22
rect 1546 18 1553 20
rect 1546 11 1551 18
rect 1568 18 1574 20
rect 1576 29 1584 31
rect 1576 27 1579 29
rect 1581 27 1584 29
rect 1576 22 1584 27
rect 1576 20 1579 22
rect 1581 20 1584 22
rect 1576 18 1584 20
rect 1586 22 1593 31
rect 1586 20 1589 22
rect 1591 20 1593 22
rect 1586 18 1593 20
rect 1608 11 1613 32
rect 1615 22 1629 38
rect 1615 20 1618 22
rect 1620 20 1629 22
rect 1631 36 1639 38
rect 1631 34 1634 36
rect 1636 34 1639 36
rect 1631 29 1639 34
rect 1631 27 1634 29
rect 1636 27 1639 29
rect 1631 20 1639 27
rect 1641 29 1649 38
rect 1641 27 1644 29
rect 1646 27 1649 29
rect 1641 20 1649 27
rect 1615 15 1627 20
rect 1615 13 1618 15
rect 1620 13 1627 15
rect 1615 11 1627 13
rect 1644 11 1649 20
rect 1651 23 1656 38
rect 1662 36 1669 38
rect 1662 34 1664 36
rect 1666 34 1669 36
rect 1662 29 1669 34
rect 1662 27 1664 29
rect 1666 27 1669 29
rect 1662 25 1669 27
rect 1651 21 1658 23
rect 1651 19 1654 21
rect 1656 19 1658 21
rect 1664 20 1669 25
rect 1671 31 1677 38
rect 1711 36 1718 38
rect 1711 34 1713 36
rect 1715 34 1718 36
rect 1711 32 1718 34
rect 1671 24 1679 31
rect 1671 22 1674 24
rect 1676 22 1679 24
rect 1671 20 1679 22
rect 1651 17 1658 19
rect 1651 11 1656 17
rect 1673 18 1679 20
rect 1681 29 1689 31
rect 1681 27 1684 29
rect 1686 27 1689 29
rect 1681 22 1689 27
rect 1681 20 1684 22
rect 1686 20 1689 22
rect 1681 18 1689 20
rect 1691 22 1698 31
rect 1691 20 1694 22
rect 1696 20 1698 22
rect 1691 18 1698 20
rect 1713 11 1718 32
rect 1720 22 1734 38
rect 1720 20 1723 22
rect 1725 20 1734 22
rect 1736 36 1744 38
rect 1736 34 1739 36
rect 1741 34 1744 36
rect 1736 29 1744 34
rect 1736 27 1739 29
rect 1741 27 1744 29
rect 1736 20 1744 27
rect 1746 29 1754 38
rect 1746 27 1749 29
rect 1751 27 1754 29
rect 1746 20 1754 27
rect 1720 15 1732 20
rect 1720 13 1723 15
rect 1725 13 1732 15
rect 1720 11 1732 13
rect 1749 11 1754 20
rect 1756 23 1761 38
rect 1769 34 1774 39
rect 1767 32 1774 34
rect 1767 30 1769 32
rect 1771 30 1774 32
rect 1767 25 1774 30
rect 1767 23 1769 25
rect 1771 23 1774 25
rect 1756 21 1763 23
rect 1767 21 1774 23
rect 1776 32 1784 39
rect 1807 36 1814 38
rect 1807 34 1809 36
rect 1811 34 1814 36
rect 1776 21 1787 32
rect 1756 19 1759 21
rect 1761 19 1763 21
rect 1756 17 1763 19
rect 1756 11 1761 17
rect 1778 15 1787 21
rect 1778 13 1780 15
rect 1782 13 1787 15
rect 1778 11 1787 13
rect 1789 11 1794 32
rect 1796 24 1801 32
rect 1807 29 1814 34
rect 1807 27 1809 29
rect 1811 27 1814 29
rect 1807 25 1814 27
rect 1796 22 1803 24
rect 1796 20 1799 22
rect 1801 20 1803 22
rect 1809 20 1814 25
rect 1816 31 1822 38
rect 1856 36 1863 38
rect 1856 34 1858 36
rect 1860 34 1863 36
rect 1856 32 1863 34
rect 1816 24 1824 31
rect 1816 22 1819 24
rect 1821 22 1824 24
rect 1816 20 1824 22
rect 1796 18 1803 20
rect 1796 11 1801 18
rect 1818 18 1824 20
rect 1826 29 1834 31
rect 1826 27 1829 29
rect 1831 27 1834 29
rect 1826 22 1834 27
rect 1826 20 1829 22
rect 1831 20 1834 22
rect 1826 18 1834 20
rect 1836 22 1843 31
rect 1836 20 1839 22
rect 1841 20 1843 22
rect 1836 18 1843 20
rect 1858 11 1863 32
rect 1865 22 1879 38
rect 1865 20 1868 22
rect 1870 20 1879 22
rect 1881 36 1889 38
rect 1881 34 1884 36
rect 1886 34 1889 36
rect 1881 29 1889 34
rect 1881 27 1884 29
rect 1886 27 1889 29
rect 1881 20 1889 27
rect 1891 29 1899 38
rect 1891 27 1894 29
rect 1896 27 1899 29
rect 1891 20 1899 27
rect 1865 15 1877 20
rect 1865 13 1868 15
rect 1870 13 1877 15
rect 1865 11 1877 13
rect 1894 11 1899 20
rect 1901 23 1906 38
rect 1912 36 1919 38
rect 1912 34 1914 36
rect 1916 34 1919 36
rect 1912 29 1919 34
rect 1912 27 1914 29
rect 1916 27 1919 29
rect 1912 25 1919 27
rect 1901 21 1908 23
rect 1901 19 1904 21
rect 1906 19 1908 21
rect 1914 20 1919 25
rect 1921 31 1927 38
rect 1961 36 1968 38
rect 1961 34 1963 36
rect 1965 34 1968 36
rect 1961 32 1968 34
rect 1921 24 1929 31
rect 1921 22 1924 24
rect 1926 22 1929 24
rect 1921 20 1929 22
rect 1901 17 1908 19
rect 1901 11 1906 17
rect 1923 18 1929 20
rect 1931 29 1939 31
rect 1931 27 1934 29
rect 1936 27 1939 29
rect 1931 22 1939 27
rect 1931 20 1934 22
rect 1936 20 1939 22
rect 1931 18 1939 20
rect 1941 22 1948 31
rect 1941 20 1944 22
rect 1946 20 1948 22
rect 1941 18 1948 20
rect 1963 11 1968 32
rect 1970 22 1984 38
rect 1970 20 1973 22
rect 1975 20 1984 22
rect 1986 36 1994 38
rect 1986 34 1989 36
rect 1991 34 1994 36
rect 1986 29 1994 34
rect 1986 27 1989 29
rect 1991 27 1994 29
rect 1986 20 1994 27
rect 1996 29 2004 38
rect 1996 27 1999 29
rect 2001 27 2004 29
rect 1996 20 2004 27
rect 1970 15 1982 20
rect 1970 13 1973 15
rect 1975 13 1982 15
rect 1970 11 1982 13
rect 1999 11 2004 20
rect 2006 23 2011 38
rect 2006 21 2013 23
rect 2006 19 2009 21
rect 2011 19 2013 21
rect 2006 17 2013 19
rect 2006 11 2011 17
<< alu1 >>
rect 33 231 1985 232
rect 23 226 2011 231
rect 23 224 54 226
rect 56 224 64 226
rect 66 224 94 226
rect 96 224 104 226
rect 106 224 122 226
rect 124 224 175 226
rect 177 224 206 226
rect 208 224 216 226
rect 218 225 1844 226
rect 218 224 366 225
rect 23 223 366 224
rect 368 223 376 225
rect 378 223 424 225
rect 426 223 434 225
rect 436 223 446 225
rect 448 223 456 225
rect 458 223 487 225
rect 489 223 540 225
rect 542 223 571 225
rect 573 223 581 225
rect 583 223 629 225
rect 631 223 639 225
rect 641 223 651 225
rect 653 223 661 225
rect 663 223 692 225
rect 694 223 745 225
rect 747 224 1844 225
rect 1846 224 1854 226
rect 1856 224 1884 226
rect 1886 224 1894 226
rect 1896 224 1912 226
rect 1914 224 1965 226
rect 1967 224 1996 226
rect 1998 224 2006 226
rect 2008 224 2011 226
rect 747 223 2011 224
rect 40 201 45 210
rect 57 214 69 218
rect 57 212 65 214
rect 67 212 69 214
rect 65 209 69 212
rect 40 200 54 201
rect 40 198 48 200
rect 50 198 51 200
rect 53 198 54 200
rect 40 197 54 198
rect 33 192 46 193
rect 33 190 38 192
rect 40 190 46 192
rect 33 189 46 190
rect 33 184 37 189
rect 65 207 66 209
rect 68 207 69 209
rect 65 192 69 207
rect 80 201 85 210
rect 97 214 109 218
rect 353 222 753 223
rect 97 212 105 214
rect 107 212 109 214
rect 80 200 94 201
rect 80 198 88 200
rect 90 198 91 200
rect 93 198 94 200
rect 80 197 94 198
rect 33 182 34 184
rect 36 182 37 184
rect 33 180 37 182
rect 64 190 69 192
rect 64 188 65 190
rect 67 188 69 190
rect 64 183 69 188
rect 64 181 65 183
rect 67 181 69 183
rect 64 179 69 181
rect 73 192 86 193
rect 73 190 78 192
rect 80 190 86 192
rect 73 189 86 190
rect 73 185 77 189
rect 105 192 109 212
rect 73 183 74 185
rect 76 183 77 185
rect 73 180 77 183
rect 104 190 109 192
rect 104 188 105 190
rect 107 188 109 190
rect 104 186 109 188
rect 104 184 105 186
rect 107 184 109 186
rect 104 183 109 184
rect 104 181 105 183
rect 107 181 109 183
rect 104 179 109 181
rect 120 216 144 217
rect 120 214 140 216
rect 142 214 144 216
rect 120 213 144 214
rect 120 194 124 213
rect 159 209 172 210
rect 159 207 167 209
rect 169 207 172 209
rect 159 205 172 207
rect 159 203 160 205
rect 162 204 172 205
rect 162 203 164 204
rect 120 192 121 194
rect 123 192 124 194
rect 120 185 124 192
rect 120 183 136 185
rect 120 181 132 183
rect 134 181 136 183
rect 120 180 136 181
rect 159 196 164 203
rect 192 209 197 210
rect 192 207 194 209
rect 196 207 197 209
rect 192 201 197 207
rect 209 214 221 218
rect 209 212 217 214
rect 219 212 221 214
rect 192 200 206 201
rect 192 198 200 200
rect 202 198 206 200
rect 192 197 206 198
rect 175 193 180 194
rect 175 192 181 193
rect 185 192 198 193
rect 175 190 176 192
rect 178 190 190 192
rect 192 190 198 192
rect 175 189 198 190
rect 175 187 189 189
rect 175 178 180 187
rect 185 186 189 187
rect 217 197 221 212
rect 217 195 218 197
rect 220 195 221 197
rect 217 192 221 195
rect 185 184 186 186
rect 188 184 189 186
rect 185 180 189 184
rect 216 190 221 192
rect 216 188 217 190
rect 219 188 221 190
rect 216 183 221 188
rect 168 172 180 178
rect 216 181 217 183
rect 219 181 221 183
rect 216 179 221 181
rect 363 213 375 217
rect 363 211 365 213
rect 367 211 375 213
rect 363 191 367 211
rect 387 200 392 209
rect 363 189 368 191
rect 363 187 365 189
rect 367 187 368 189
rect 363 182 368 187
rect 363 180 365 182
rect 367 180 368 182
rect 378 199 392 200
rect 378 197 379 199
rect 381 197 382 199
rect 384 197 392 199
rect 378 196 392 197
rect 410 200 415 209
rect 427 213 439 217
rect 427 211 435 213
rect 437 211 439 213
rect 435 208 439 211
rect 410 199 424 200
rect 410 197 418 199
rect 420 197 421 199
rect 423 197 424 199
rect 410 196 424 197
rect 386 191 399 192
rect 386 189 392 191
rect 394 189 399 191
rect 386 188 399 189
rect 363 178 368 180
rect 32 166 221 167
rect 395 182 399 188
rect 395 180 396 182
rect 398 180 399 182
rect 395 179 399 180
rect 403 191 416 192
rect 403 189 404 191
rect 406 189 408 191
rect 410 189 416 191
rect 403 188 416 189
rect 403 179 407 188
rect 435 206 436 208
rect 438 206 439 208
rect 435 191 439 206
rect 434 189 439 191
rect 434 187 435 189
rect 437 187 439 189
rect 434 182 439 187
rect 434 180 435 182
rect 437 180 439 182
rect 434 178 439 180
rect 443 213 455 217
rect 443 211 445 213
rect 447 211 455 213
rect 520 215 544 216
rect 443 200 447 211
rect 520 213 522 215
rect 524 213 544 215
rect 520 212 544 213
rect 443 198 444 200
rect 446 198 447 200
rect 443 191 447 198
rect 467 208 472 209
rect 467 206 468 208
rect 470 206 472 208
rect 467 200 472 206
rect 443 189 448 191
rect 443 187 445 189
rect 447 187 448 189
rect 443 182 448 187
rect 443 180 445 182
rect 447 180 448 182
rect 458 199 472 200
rect 458 197 462 199
rect 464 197 472 199
rect 458 196 472 197
rect 492 208 505 209
rect 492 206 495 208
rect 497 206 505 208
rect 492 204 505 206
rect 492 203 502 204
rect 500 202 502 203
rect 504 202 505 204
rect 484 192 489 193
rect 466 191 479 192
rect 483 191 489 192
rect 466 189 472 191
rect 474 189 486 191
rect 488 189 489 191
rect 466 188 489 189
rect 475 186 489 188
rect 500 195 505 202
rect 443 178 448 180
rect 475 179 479 186
rect 484 177 489 186
rect 484 175 496 177
rect 484 173 492 175
rect 494 173 496 175
rect 484 171 496 173
rect 540 184 544 212
rect 528 182 544 184
rect 528 180 530 182
rect 532 180 544 182
rect 528 179 544 180
rect 568 213 580 217
rect 568 211 570 213
rect 572 211 580 213
rect 568 191 572 211
rect 592 200 597 209
rect 568 189 573 191
rect 568 187 570 189
rect 572 187 573 189
rect 568 186 573 187
rect 568 184 570 186
rect 572 184 573 186
rect 568 182 573 184
rect 568 180 570 182
rect 572 180 573 182
rect 583 199 597 200
rect 583 197 584 199
rect 586 197 587 199
rect 589 197 597 199
rect 583 196 597 197
rect 615 200 620 209
rect 632 213 644 217
rect 632 211 640 213
rect 642 211 644 213
rect 640 208 644 211
rect 615 199 629 200
rect 615 197 623 199
rect 625 197 626 199
rect 628 197 629 199
rect 615 196 629 197
rect 591 191 604 192
rect 591 189 597 191
rect 599 189 604 191
rect 591 188 604 189
rect 568 178 573 180
rect 600 182 604 188
rect 600 180 601 182
rect 603 180 604 182
rect 600 179 604 180
rect 608 191 621 192
rect 608 189 609 191
rect 611 189 613 191
rect 615 189 621 191
rect 608 188 621 189
rect 608 179 612 188
rect 640 206 641 208
rect 643 206 644 208
rect 640 191 644 206
rect 639 189 644 191
rect 639 187 640 189
rect 642 187 644 189
rect 639 182 644 187
rect 639 180 640 182
rect 642 180 644 182
rect 639 178 644 180
rect 648 213 660 217
rect 648 211 650 213
rect 652 211 660 213
rect 725 215 749 216
rect 648 198 652 211
rect 725 213 727 215
rect 729 213 749 215
rect 725 212 749 213
rect 648 196 649 198
rect 651 196 652 198
rect 648 191 652 196
rect 672 208 677 209
rect 672 206 673 208
rect 675 206 677 208
rect 672 200 677 206
rect 648 189 653 191
rect 648 187 650 189
rect 652 187 653 189
rect 648 182 653 187
rect 648 180 650 182
rect 652 180 653 182
rect 663 199 677 200
rect 663 197 667 199
rect 669 197 677 199
rect 663 196 677 197
rect 697 208 710 209
rect 697 206 700 208
rect 702 206 710 208
rect 697 204 710 206
rect 697 203 707 204
rect 705 202 707 203
rect 709 202 710 204
rect 689 192 694 193
rect 671 191 684 192
rect 688 191 694 192
rect 671 189 677 191
rect 679 189 691 191
rect 693 189 694 191
rect 671 188 694 189
rect 680 186 694 188
rect 705 195 710 202
rect 648 178 653 180
rect 680 179 684 186
rect 689 177 694 186
rect 689 175 701 177
rect 689 173 697 175
rect 699 173 701 175
rect 689 171 701 173
rect 745 184 749 212
rect 1830 201 1835 210
rect 1847 214 1859 218
rect 1847 212 1855 214
rect 1857 212 1859 214
rect 1855 209 1859 212
rect 1830 200 1844 201
rect 1830 198 1838 200
rect 1840 198 1841 200
rect 1843 198 1844 200
rect 1830 197 1844 198
rect 733 182 749 184
rect 733 180 735 182
rect 737 180 746 182
rect 748 180 749 182
rect 1823 192 1836 193
rect 1823 190 1828 192
rect 1830 190 1836 192
rect 1823 189 1836 190
rect 1823 184 1827 189
rect 1855 207 1856 209
rect 1858 207 1859 209
rect 1855 192 1859 207
rect 1870 201 1875 210
rect 1887 214 1899 218
rect 1887 212 1895 214
rect 1897 212 1899 214
rect 1870 200 1884 201
rect 1870 198 1878 200
rect 1880 198 1881 200
rect 1883 198 1884 200
rect 1870 197 1884 198
rect 1823 182 1824 184
rect 1826 182 1827 184
rect 1823 180 1827 182
rect 1854 190 1859 192
rect 1854 188 1855 190
rect 1857 188 1859 190
rect 1854 183 1859 188
rect 733 179 749 180
rect 1854 181 1855 183
rect 1857 181 1859 183
rect 1854 179 1859 181
rect 1863 192 1876 193
rect 1863 190 1868 192
rect 1870 190 1876 192
rect 1863 189 1876 190
rect 1863 185 1867 189
rect 1895 192 1899 212
rect 1863 183 1864 185
rect 1866 183 1867 185
rect 1863 180 1867 183
rect 1894 190 1899 192
rect 1894 188 1895 190
rect 1897 188 1899 190
rect 1894 186 1899 188
rect 1894 184 1895 186
rect 1897 184 1899 186
rect 1894 183 1899 184
rect 1894 181 1895 183
rect 1897 181 1899 183
rect 1894 179 1899 181
rect 1910 216 1934 217
rect 1910 214 1930 216
rect 1932 214 1934 216
rect 1910 213 1934 214
rect 1910 185 1914 213
rect 1949 209 1962 210
rect 1949 207 1957 209
rect 1959 207 1962 209
rect 1949 205 1962 207
rect 1949 203 1950 205
rect 1952 204 1962 205
rect 1952 203 1954 204
rect 1910 183 1926 185
rect 1910 181 1922 183
rect 1924 181 1926 183
rect 1910 180 1926 181
rect 1949 196 1954 203
rect 1982 209 1987 210
rect 1982 207 1984 209
rect 1986 207 1987 209
rect 1982 201 1987 207
rect 1999 214 2011 218
rect 1999 212 2007 214
rect 2009 212 2011 214
rect 1982 200 1996 201
rect 1982 198 1990 200
rect 1992 198 1996 200
rect 1982 197 1996 198
rect 1965 193 1970 194
rect 1965 192 1971 193
rect 1975 192 1988 193
rect 1965 190 1966 192
rect 1968 190 1980 192
rect 1982 190 1988 192
rect 1965 189 1988 190
rect 1965 187 1979 189
rect 1965 178 1970 187
rect 1975 186 1979 187
rect 2007 197 2011 212
rect 2007 195 2008 197
rect 2010 195 2011 197
rect 2007 192 2011 195
rect 1975 184 1976 186
rect 1978 184 1979 186
rect 1975 180 1979 184
rect 2006 190 2011 192
rect 2006 188 2007 190
rect 2009 188 2011 190
rect 2006 183 2011 188
rect 1958 172 1970 178
rect 2006 181 2007 183
rect 2009 181 2011 183
rect 2006 179 2011 181
rect 1822 166 2011 167
rect 32 164 64 166
rect 66 164 104 166
rect 106 164 142 166
rect 144 164 216 166
rect 218 164 221 166
rect 32 159 221 164
rect 362 165 756 166
rect 362 163 366 165
rect 368 163 434 165
rect 436 163 446 165
rect 448 163 520 165
rect 522 163 571 165
rect 573 163 639 165
rect 641 163 651 165
rect 653 163 725 165
rect 727 163 756 165
rect 362 159 756 163
rect 1822 164 1854 166
rect 1856 164 1894 166
rect 1896 164 1932 166
rect 1934 164 2006 166
rect 2008 164 2011 166
rect 32 158 1775 159
rect 1822 158 2011 164
rect 32 154 2011 158
rect 32 152 36 154
rect 38 152 104 154
rect 106 152 116 154
rect 118 152 190 154
rect 192 152 240 154
rect 242 152 314 154
rect 316 153 778 154
rect 316 152 394 153
rect 32 151 394 152
rect 396 151 434 153
rect 436 151 472 153
rect 474 151 546 153
rect 548 151 599 153
rect 601 151 639 153
rect 641 151 677 153
rect 679 151 751 153
rect 753 152 778 153
rect 780 152 818 154
rect 820 152 892 154
rect 894 152 923 154
rect 925 152 997 154
rect 999 152 1028 154
rect 1030 152 1068 154
rect 1070 152 1142 154
rect 1144 152 1173 154
rect 1175 152 1247 154
rect 1249 152 1278 154
rect 1280 152 1318 154
rect 1320 152 1392 154
rect 1394 152 1423 154
rect 1425 152 1497 154
rect 1499 152 1528 154
rect 1530 152 1568 154
rect 1570 152 1642 154
rect 1644 152 1673 154
rect 1675 152 1747 154
rect 1749 152 1826 154
rect 1828 152 1894 154
rect 1896 152 1906 154
rect 1908 152 1980 154
rect 1982 152 2011 154
rect 753 151 2011 152
rect 33 137 38 139
rect 33 135 35 137
rect 37 135 38 137
rect 33 130 38 135
rect 33 128 35 130
rect 37 128 38 130
rect 33 126 38 128
rect 65 137 69 138
rect 65 135 66 137
rect 68 135 69 137
rect 33 122 37 126
rect 33 121 38 122
rect 33 119 35 121
rect 37 119 38 121
rect 33 115 38 119
rect 65 129 69 135
rect 56 128 69 129
rect 56 126 62 128
rect 64 126 69 128
rect 56 125 69 126
rect 73 129 77 138
rect 104 137 109 139
rect 73 128 86 129
rect 73 126 74 128
rect 76 126 78 128
rect 80 126 86 128
rect 73 125 86 126
rect 33 106 37 115
rect 48 120 62 121
rect 48 118 49 120
rect 51 118 52 120
rect 54 118 62 120
rect 48 117 62 118
rect 33 104 35 106
rect 37 104 45 106
rect 33 100 45 104
rect 57 108 62 117
rect 80 120 94 121
rect 80 118 88 120
rect 90 118 91 120
rect 93 118 94 120
rect 80 117 94 118
rect 104 135 105 137
rect 107 135 109 137
rect 104 130 109 135
rect 104 128 105 130
rect 107 128 109 130
rect 104 126 109 128
rect 80 108 85 117
rect 105 111 109 126
rect 105 109 106 111
rect 108 109 109 111
rect 105 106 109 109
rect 97 104 105 106
rect 107 104 109 106
rect 97 100 109 104
rect 113 137 118 139
rect 113 135 115 137
rect 117 135 118 137
rect 154 144 166 146
rect 154 142 162 144
rect 164 142 166 144
rect 154 140 166 142
rect 113 130 118 135
rect 113 128 115 130
rect 117 128 118 130
rect 113 126 118 128
rect 113 119 117 126
rect 113 117 114 119
rect 116 117 117 119
rect 113 106 117 117
rect 145 131 149 138
rect 154 131 159 140
rect 145 129 159 131
rect 136 128 159 129
rect 136 126 142 128
rect 144 126 156 128
rect 158 126 159 128
rect 136 125 149 126
rect 153 125 159 126
rect 154 124 159 125
rect 128 120 142 121
rect 128 118 132 120
rect 134 118 142 120
rect 128 117 142 118
rect 113 104 115 106
rect 117 104 125 106
rect 113 100 125 104
rect 137 111 142 117
rect 137 109 138 111
rect 140 109 142 111
rect 137 108 142 109
rect 170 115 175 122
rect 198 137 214 138
rect 198 135 200 137
rect 202 135 214 137
rect 198 133 214 135
rect 170 114 172 115
rect 162 113 172 114
rect 174 113 175 115
rect 162 111 175 113
rect 162 109 165 111
rect 167 109 175 111
rect 162 108 175 109
rect 210 110 214 133
rect 210 108 211 110
rect 213 108 214 110
rect 210 105 214 108
rect 190 104 214 105
rect 190 102 192 104
rect 194 102 214 104
rect 190 101 214 102
rect 237 137 242 139
rect 237 135 239 137
rect 241 135 242 137
rect 362 150 781 151
rect 278 140 290 146
rect 237 130 242 135
rect 237 128 239 130
rect 241 128 242 130
rect 237 126 242 128
rect 237 109 241 126
rect 269 131 273 138
rect 278 131 283 140
rect 269 129 283 131
rect 260 128 283 129
rect 260 126 266 128
rect 268 126 280 128
rect 282 126 283 128
rect 260 125 273 126
rect 277 125 283 126
rect 278 124 283 125
rect 252 120 266 121
rect 252 118 256 120
rect 258 118 266 120
rect 252 117 266 118
rect 237 107 238 109
rect 240 107 241 109
rect 237 106 241 107
rect 237 104 239 106
rect 241 104 249 106
rect 237 100 249 104
rect 261 111 266 117
rect 261 109 262 111
rect 264 109 266 111
rect 261 108 266 109
rect 294 115 299 122
rect 322 137 338 138
rect 322 135 324 137
rect 326 135 338 137
rect 322 133 338 135
rect 294 114 296 115
rect 286 113 296 114
rect 298 113 299 115
rect 286 111 299 113
rect 286 109 289 111
rect 291 109 299 111
rect 286 108 299 109
rect 334 105 338 133
rect 363 135 367 137
rect 363 133 364 135
rect 366 133 367 135
rect 363 128 367 133
rect 394 136 399 138
rect 363 127 376 128
rect 363 125 368 127
rect 370 125 376 127
rect 363 124 376 125
rect 370 119 384 120
rect 370 117 378 119
rect 380 117 381 119
rect 383 117 384 119
rect 370 116 384 117
rect 394 134 395 136
rect 397 134 399 136
rect 394 129 399 134
rect 394 127 395 129
rect 397 127 399 129
rect 394 125 399 127
rect 370 107 375 116
rect 395 110 399 125
rect 403 134 407 137
rect 403 132 404 134
rect 406 132 407 134
rect 403 128 407 132
rect 434 136 439 138
rect 403 127 416 128
rect 403 125 408 127
rect 410 125 416 127
rect 403 124 416 125
rect 395 108 396 110
rect 398 108 399 110
rect 314 104 338 105
rect 395 105 399 108
rect 410 119 424 120
rect 410 117 418 119
rect 420 117 421 119
rect 423 117 424 119
rect 410 116 424 117
rect 434 134 435 136
rect 437 134 439 136
rect 434 133 439 134
rect 434 131 435 133
rect 437 131 439 133
rect 434 129 439 131
rect 434 127 435 129
rect 437 127 439 129
rect 434 125 439 127
rect 410 107 415 116
rect 314 102 316 104
rect 318 102 335 104
rect 337 102 338 104
rect 314 101 338 102
rect 387 103 395 105
rect 397 103 399 105
rect 435 105 439 125
rect 387 99 399 103
rect 427 103 435 105
rect 437 103 439 105
rect 427 99 439 103
rect 450 136 466 137
rect 450 134 462 136
rect 464 134 466 136
rect 450 132 466 134
rect 450 104 454 132
rect 498 139 510 145
rect 505 130 510 139
rect 515 133 519 137
rect 515 131 516 133
rect 518 131 519 133
rect 546 136 551 138
rect 515 130 519 131
rect 489 114 494 121
rect 505 128 519 130
rect 505 127 528 128
rect 505 125 506 127
rect 508 125 520 127
rect 522 125 528 127
rect 505 124 511 125
rect 515 124 528 125
rect 505 123 510 124
rect 489 112 490 114
rect 492 113 494 114
rect 492 112 502 113
rect 489 110 502 112
rect 489 108 497 110
rect 499 108 502 110
rect 489 107 502 108
rect 522 119 536 120
rect 522 117 530 119
rect 532 117 536 119
rect 522 116 536 117
rect 546 134 547 136
rect 549 134 551 136
rect 546 129 551 134
rect 546 127 547 129
rect 549 127 551 129
rect 546 125 551 127
rect 522 110 527 116
rect 522 108 524 110
rect 526 108 527 110
rect 522 107 527 108
rect 547 122 551 125
rect 568 135 572 137
rect 568 133 569 135
rect 571 133 572 135
rect 568 128 572 133
rect 599 136 604 138
rect 568 127 581 128
rect 568 125 573 127
rect 575 125 581 127
rect 568 124 581 125
rect 547 120 548 122
rect 550 120 551 122
rect 450 103 474 104
rect 450 101 470 103
rect 472 101 474 103
rect 547 105 551 120
rect 575 119 589 120
rect 575 117 583 119
rect 585 117 586 119
rect 588 117 589 119
rect 575 116 589 117
rect 599 134 600 136
rect 602 134 604 136
rect 599 129 604 134
rect 599 127 600 129
rect 602 127 604 129
rect 599 125 604 127
rect 575 107 580 116
rect 600 110 604 125
rect 608 134 612 137
rect 608 132 609 134
rect 611 132 612 134
rect 608 128 612 132
rect 639 136 644 138
rect 608 127 621 128
rect 608 125 613 127
rect 615 125 621 127
rect 608 124 621 125
rect 600 108 601 110
rect 603 108 604 110
rect 450 100 474 101
rect 539 103 547 105
rect 549 103 551 105
rect 600 105 604 108
rect 615 119 629 120
rect 615 117 623 119
rect 625 117 626 119
rect 628 117 629 119
rect 615 116 629 117
rect 639 134 640 136
rect 642 134 644 136
rect 639 133 644 134
rect 639 131 640 133
rect 642 131 644 133
rect 639 129 644 131
rect 639 127 640 129
rect 642 127 644 129
rect 639 125 644 127
rect 615 107 620 116
rect 23 94 342 95
rect 539 99 551 103
rect 592 103 600 105
rect 602 103 604 105
rect 640 105 644 125
rect 592 99 604 103
rect 632 103 640 105
rect 642 103 644 105
rect 632 99 644 103
rect 655 136 671 137
rect 655 134 667 136
rect 669 134 671 136
rect 655 132 671 134
rect 655 118 659 132
rect 703 139 715 145
rect 710 130 715 139
rect 720 133 724 137
rect 720 131 721 133
rect 723 131 724 133
rect 775 141 788 145
rect 775 139 777 141
rect 751 136 756 138
rect 720 130 724 131
rect 655 116 656 118
rect 658 116 659 118
rect 655 104 659 116
rect 694 114 699 121
rect 710 128 724 130
rect 710 127 733 128
rect 710 125 711 127
rect 713 125 725 127
rect 727 125 733 127
rect 710 124 716 125
rect 720 124 733 125
rect 710 123 715 124
rect 694 112 695 114
rect 697 113 699 114
rect 697 112 707 113
rect 694 110 707 112
rect 694 108 702 110
rect 704 108 707 110
rect 694 107 707 108
rect 727 119 741 120
rect 727 117 735 119
rect 737 117 741 119
rect 727 116 741 117
rect 751 134 752 136
rect 754 134 756 136
rect 751 129 756 134
rect 751 127 752 129
rect 754 127 756 129
rect 751 125 756 127
rect 727 110 732 116
rect 727 108 729 110
rect 731 108 732 110
rect 727 107 732 108
rect 752 122 756 125
rect 752 120 753 122
rect 755 120 756 122
rect 655 103 679 104
rect 655 101 675 103
rect 677 101 679 103
rect 752 105 756 120
rect 775 134 779 139
rect 775 132 777 134
rect 775 113 779 132
rect 807 137 811 138
rect 807 135 808 137
rect 810 135 811 137
rect 807 129 811 135
rect 790 127 811 129
rect 790 125 804 127
rect 806 125 811 127
rect 815 137 820 139
rect 815 135 817 137
rect 819 135 820 137
rect 856 140 868 146
rect 815 130 820 135
rect 815 128 817 130
rect 819 128 820 130
rect 815 126 820 128
rect 815 121 819 126
rect 775 111 780 113
rect 775 109 777 111
rect 779 109 780 111
rect 775 107 780 109
rect 790 120 819 121
rect 790 118 794 120
rect 796 118 819 120
rect 790 117 819 118
rect 807 108 811 117
rect 655 100 679 101
rect 744 103 752 105
rect 754 103 756 105
rect 744 99 756 103
rect 815 106 819 117
rect 847 131 851 138
rect 856 131 861 140
rect 847 129 861 131
rect 838 128 861 129
rect 838 126 844 128
rect 846 126 858 128
rect 860 126 861 128
rect 838 125 851 126
rect 855 125 861 126
rect 856 124 861 125
rect 830 120 844 121
rect 830 118 834 120
rect 836 118 844 120
rect 830 117 844 118
rect 815 104 817 106
rect 819 104 827 106
rect 815 100 827 104
rect 839 111 844 117
rect 839 109 840 111
rect 842 109 844 111
rect 839 108 844 109
rect 872 115 877 122
rect 900 137 916 138
rect 900 135 902 137
rect 904 135 916 137
rect 900 133 916 135
rect 872 114 874 115
rect 864 113 874 114
rect 876 113 877 115
rect 864 111 877 113
rect 864 109 867 111
rect 869 109 877 111
rect 864 108 877 109
rect 912 111 916 133
rect 912 109 913 111
rect 915 109 916 111
rect 912 105 916 109
rect 892 104 916 105
rect 892 102 894 104
rect 896 102 916 104
rect 892 101 916 102
rect 920 137 925 139
rect 920 135 922 137
rect 924 135 925 137
rect 961 140 973 146
rect 1025 145 1029 146
rect 920 130 925 135
rect 920 128 922 130
rect 924 128 925 130
rect 920 126 925 128
rect 920 106 924 126
rect 952 131 956 138
rect 961 131 966 140
rect 1025 141 1038 145
rect 1025 139 1027 141
rect 952 129 966 131
rect 943 128 955 129
rect 943 126 949 128
rect 951 127 955 128
rect 957 128 966 129
rect 957 127 963 128
rect 951 126 963 127
rect 965 126 966 128
rect 943 125 956 126
rect 960 125 966 126
rect 961 124 966 125
rect 935 120 949 121
rect 935 118 939 120
rect 941 118 949 120
rect 935 117 949 118
rect 920 104 922 106
rect 924 104 932 106
rect 920 100 932 104
rect 944 111 949 117
rect 944 109 945 111
rect 947 109 949 111
rect 944 108 949 109
rect 977 115 982 122
rect 1005 137 1021 138
rect 1005 135 1007 137
rect 1009 135 1021 137
rect 1005 133 1021 135
rect 977 114 979 115
rect 969 113 979 114
rect 981 113 982 115
rect 969 111 982 113
rect 969 109 972 111
rect 974 109 982 111
rect 969 108 982 109
rect 1017 105 1021 133
rect 1025 134 1029 139
rect 1025 132 1027 134
rect 1025 129 1029 132
rect 1057 137 1061 138
rect 1057 135 1058 137
rect 1060 135 1061 137
rect 1025 127 1026 129
rect 1028 127 1029 129
rect 1025 113 1029 127
rect 1057 129 1061 135
rect 1040 127 1061 129
rect 1040 125 1054 127
rect 1056 125 1061 127
rect 1065 137 1070 139
rect 1065 135 1067 137
rect 1069 135 1070 137
rect 1106 140 1118 146
rect 1065 130 1070 135
rect 1065 128 1067 130
rect 1069 128 1070 130
rect 1065 126 1070 128
rect 1065 121 1069 126
rect 1025 111 1030 113
rect 1025 109 1027 111
rect 1029 109 1030 111
rect 1025 107 1030 109
rect 1040 120 1069 121
rect 1040 118 1044 120
rect 1046 118 1069 120
rect 1040 117 1069 118
rect 1057 108 1061 117
rect 997 104 1021 105
rect 997 102 999 104
rect 1001 102 1018 104
rect 1020 102 1021 104
rect 997 101 1021 102
rect 1065 106 1069 117
rect 1097 131 1101 138
rect 1106 131 1111 140
rect 1097 129 1111 131
rect 1088 128 1111 129
rect 1088 126 1094 128
rect 1096 126 1108 128
rect 1110 126 1111 128
rect 1088 125 1101 126
rect 1105 125 1111 126
rect 1106 124 1111 125
rect 1080 120 1094 121
rect 1080 118 1084 120
rect 1086 118 1094 120
rect 1080 117 1094 118
rect 1065 104 1067 106
rect 1069 104 1077 106
rect 1065 100 1077 104
rect 1089 111 1094 117
rect 1089 109 1090 111
rect 1092 109 1094 111
rect 1089 108 1094 109
rect 1122 115 1127 122
rect 1150 137 1166 138
rect 1150 135 1152 137
rect 1154 135 1166 137
rect 1150 133 1166 135
rect 1122 114 1124 115
rect 1114 113 1124 114
rect 1126 113 1127 115
rect 1114 111 1127 113
rect 1114 109 1117 111
rect 1119 109 1127 111
rect 1114 108 1127 109
rect 1162 111 1166 133
rect 1162 109 1163 111
rect 1165 109 1166 111
rect 1162 105 1166 109
rect 1142 104 1166 105
rect 1142 102 1144 104
rect 1146 102 1166 104
rect 1142 101 1166 102
rect 1170 137 1175 139
rect 1170 135 1172 137
rect 1174 135 1175 137
rect 1211 140 1223 146
rect 1275 145 1279 146
rect 1170 130 1175 135
rect 1170 128 1172 130
rect 1174 128 1175 130
rect 1170 126 1175 128
rect 1170 106 1174 126
rect 1202 131 1206 138
rect 1211 131 1216 140
rect 1275 141 1288 145
rect 1275 139 1277 141
rect 1202 129 1216 131
rect 1193 128 1207 129
rect 1193 126 1199 128
rect 1201 127 1207 128
rect 1209 128 1216 129
rect 1209 127 1213 128
rect 1201 126 1213 127
rect 1215 126 1216 128
rect 1193 125 1206 126
rect 1210 125 1216 126
rect 1211 124 1216 125
rect 1185 120 1199 121
rect 1185 118 1189 120
rect 1191 118 1199 120
rect 1185 117 1199 118
rect 1170 104 1172 106
rect 1174 104 1182 106
rect 1170 100 1182 104
rect 1194 111 1199 117
rect 1194 109 1195 111
rect 1197 109 1199 111
rect 1194 108 1199 109
rect 1227 115 1232 122
rect 1255 137 1271 138
rect 1255 135 1257 137
rect 1259 135 1271 137
rect 1255 133 1271 135
rect 1227 114 1229 115
rect 1219 113 1229 114
rect 1231 113 1232 115
rect 1219 111 1232 113
rect 1219 109 1222 111
rect 1224 109 1232 111
rect 1219 108 1232 109
rect 1267 105 1271 133
rect 1275 134 1279 139
rect 1275 132 1277 134
rect 1275 129 1279 132
rect 1307 137 1311 138
rect 1307 135 1308 137
rect 1310 135 1311 137
rect 1275 127 1276 129
rect 1278 127 1279 129
rect 1275 113 1279 127
rect 1307 129 1311 135
rect 1290 127 1311 129
rect 1290 125 1304 127
rect 1306 125 1311 127
rect 1315 137 1320 139
rect 1315 135 1317 137
rect 1319 135 1320 137
rect 1356 140 1368 146
rect 1315 130 1320 135
rect 1315 128 1317 130
rect 1319 128 1320 130
rect 1315 126 1320 128
rect 1315 121 1319 126
rect 1275 111 1280 113
rect 1275 109 1277 111
rect 1279 109 1280 111
rect 1275 107 1280 109
rect 1290 120 1319 121
rect 1290 118 1294 120
rect 1296 118 1319 120
rect 1290 117 1319 118
rect 1307 108 1311 117
rect 1247 104 1268 105
rect 1247 102 1249 104
rect 1251 103 1268 104
rect 1270 103 1271 105
rect 1251 102 1271 103
rect 1247 101 1271 102
rect 1315 106 1319 117
rect 1347 131 1351 138
rect 1356 131 1361 140
rect 1347 129 1361 131
rect 1338 128 1361 129
rect 1338 126 1344 128
rect 1346 126 1358 128
rect 1360 126 1361 128
rect 1338 125 1351 126
rect 1355 125 1361 126
rect 1356 124 1361 125
rect 1330 120 1344 121
rect 1330 118 1334 120
rect 1336 118 1344 120
rect 1330 117 1344 118
rect 1315 104 1317 106
rect 1319 104 1327 106
rect 1315 100 1327 104
rect 1339 111 1344 117
rect 1339 109 1340 111
rect 1342 109 1344 111
rect 1339 108 1344 109
rect 1372 115 1377 122
rect 1400 137 1416 138
rect 1400 135 1402 137
rect 1404 135 1416 137
rect 1400 133 1416 135
rect 1372 114 1374 115
rect 1364 113 1374 114
rect 1376 113 1377 115
rect 1364 111 1377 113
rect 1364 109 1367 111
rect 1369 109 1377 111
rect 1364 108 1377 109
rect 1412 111 1416 133
rect 1412 109 1413 111
rect 1415 109 1416 111
rect 1412 105 1416 109
rect 1392 104 1416 105
rect 1392 102 1394 104
rect 1396 102 1416 104
rect 1392 101 1416 102
rect 1420 137 1425 139
rect 1420 135 1422 137
rect 1424 135 1425 137
rect 1461 140 1473 146
rect 1525 145 1529 146
rect 1420 130 1425 135
rect 1420 128 1422 130
rect 1424 128 1425 130
rect 1420 126 1425 128
rect 1420 106 1424 126
rect 1452 131 1456 138
rect 1461 131 1466 140
rect 1525 141 1538 145
rect 1525 139 1527 141
rect 1452 129 1466 131
rect 1443 128 1457 129
rect 1443 126 1449 128
rect 1451 127 1457 128
rect 1459 128 1466 129
rect 1459 127 1463 128
rect 1451 126 1463 127
rect 1465 126 1466 128
rect 1443 125 1456 126
rect 1460 125 1466 126
rect 1461 124 1466 125
rect 1435 120 1449 121
rect 1435 118 1439 120
rect 1441 118 1449 120
rect 1435 117 1449 118
rect 1420 104 1422 106
rect 1424 104 1432 106
rect 1420 100 1432 104
rect 1444 111 1449 117
rect 1444 109 1445 111
rect 1447 109 1449 111
rect 1444 108 1449 109
rect 1477 115 1482 122
rect 1505 137 1521 138
rect 1505 135 1507 137
rect 1509 135 1521 137
rect 1505 133 1521 135
rect 1477 114 1479 115
rect 1469 113 1479 114
rect 1481 113 1482 115
rect 1469 111 1482 113
rect 1469 109 1472 111
rect 1474 109 1482 111
rect 1469 108 1482 109
rect 1517 105 1521 133
rect 1525 134 1529 139
rect 1525 132 1527 134
rect 1525 129 1529 132
rect 1557 137 1561 138
rect 1557 135 1558 137
rect 1560 135 1561 137
rect 1525 127 1526 129
rect 1528 127 1529 129
rect 1525 113 1529 127
rect 1557 129 1561 135
rect 1540 127 1561 129
rect 1540 125 1554 127
rect 1556 125 1561 127
rect 1565 137 1570 139
rect 1565 135 1567 137
rect 1569 135 1570 137
rect 1606 140 1618 146
rect 1565 130 1570 135
rect 1565 128 1567 130
rect 1569 128 1570 130
rect 1565 126 1570 128
rect 1565 121 1569 126
rect 1525 111 1530 113
rect 1525 109 1527 111
rect 1529 109 1530 111
rect 1525 107 1530 109
rect 1540 120 1569 121
rect 1540 118 1544 120
rect 1546 118 1569 120
rect 1540 117 1569 118
rect 1557 108 1561 117
rect 1497 104 1518 105
rect 1497 102 1499 104
rect 1501 103 1518 104
rect 1520 103 1521 105
rect 1501 102 1521 103
rect 1497 101 1521 102
rect 1565 106 1569 117
rect 1597 131 1601 138
rect 1606 131 1611 140
rect 1597 129 1611 131
rect 1588 128 1611 129
rect 1588 126 1594 128
rect 1596 126 1608 128
rect 1610 126 1611 128
rect 1588 125 1601 126
rect 1605 125 1611 126
rect 1606 124 1611 125
rect 1580 120 1594 121
rect 1580 118 1584 120
rect 1586 118 1594 120
rect 1580 117 1594 118
rect 1565 104 1567 106
rect 1569 104 1577 106
rect 1565 100 1577 104
rect 1589 111 1594 117
rect 1589 109 1590 111
rect 1592 109 1594 111
rect 1589 108 1594 109
rect 1622 115 1627 122
rect 1650 137 1666 138
rect 1650 135 1652 137
rect 1654 135 1666 137
rect 1650 133 1666 135
rect 1622 114 1624 115
rect 1614 113 1624 114
rect 1626 113 1627 115
rect 1614 111 1627 113
rect 1614 109 1617 111
rect 1619 109 1627 111
rect 1614 108 1627 109
rect 1662 111 1666 133
rect 1662 109 1663 111
rect 1665 109 1666 111
rect 1662 105 1666 109
rect 1642 104 1666 105
rect 1642 102 1644 104
rect 1646 102 1666 104
rect 1642 101 1666 102
rect 1670 137 1675 139
rect 1670 135 1672 137
rect 1674 135 1675 137
rect 1711 140 1723 146
rect 1670 130 1675 135
rect 1670 128 1672 130
rect 1674 128 1675 130
rect 1670 126 1675 128
rect 1670 106 1674 126
rect 1702 131 1706 138
rect 1711 131 1716 140
rect 1702 129 1716 131
rect 1693 128 1716 129
rect 1693 126 1699 128
rect 1701 126 1713 128
rect 1715 126 1716 128
rect 1693 125 1706 126
rect 1710 125 1716 126
rect 1711 124 1716 125
rect 1685 120 1699 121
rect 1685 118 1689 120
rect 1691 118 1699 120
rect 1685 117 1699 118
rect 1670 104 1672 106
rect 1674 104 1682 106
rect 1670 100 1682 104
rect 1694 111 1699 117
rect 1694 109 1695 111
rect 1697 109 1699 111
rect 1694 108 1699 109
rect 1727 115 1732 122
rect 1755 137 1771 138
rect 1755 135 1757 137
rect 1759 135 1771 137
rect 1755 133 1771 135
rect 1727 114 1729 115
rect 1719 113 1729 114
rect 1731 113 1732 115
rect 1719 111 1732 113
rect 1719 109 1722 111
rect 1724 109 1732 111
rect 1719 108 1732 109
rect 1767 105 1771 133
rect 1747 104 1771 105
rect 1747 102 1749 104
rect 1751 102 1768 104
rect 1770 102 1771 104
rect 1747 101 1771 102
rect 1823 137 1828 139
rect 1823 135 1825 137
rect 1827 135 1828 137
rect 1823 130 1828 135
rect 1823 128 1825 130
rect 1827 128 1828 130
rect 1823 126 1828 128
rect 1855 137 1859 138
rect 1855 135 1856 137
rect 1858 135 1859 137
rect 1823 106 1827 126
rect 1855 129 1859 135
rect 1846 128 1859 129
rect 1846 126 1852 128
rect 1854 126 1859 128
rect 1846 125 1859 126
rect 1863 129 1867 138
rect 1894 137 1899 139
rect 1863 128 1876 129
rect 1863 126 1864 128
rect 1866 126 1868 128
rect 1870 126 1876 128
rect 1863 125 1876 126
rect 1838 120 1852 121
rect 1838 118 1839 120
rect 1841 118 1842 120
rect 1844 118 1852 120
rect 1838 117 1852 118
rect 1823 104 1825 106
rect 1827 104 1835 106
rect 1823 100 1835 104
rect 1847 108 1852 117
rect 1870 120 1884 121
rect 1870 118 1878 120
rect 1880 118 1881 120
rect 1883 118 1884 120
rect 1870 117 1884 118
rect 1894 135 1895 137
rect 1897 135 1899 137
rect 1894 130 1899 135
rect 1894 128 1895 130
rect 1897 128 1899 130
rect 1894 126 1899 128
rect 1870 108 1875 117
rect 1895 111 1899 126
rect 1895 109 1896 111
rect 1898 109 1899 111
rect 1895 106 1899 109
rect 1887 104 1895 106
rect 1897 104 1899 106
rect 1887 100 1899 104
rect 1903 137 1908 139
rect 1903 135 1905 137
rect 1907 135 1908 137
rect 1944 144 1956 146
rect 1944 142 1952 144
rect 1954 142 1956 144
rect 1944 140 1956 142
rect 1903 130 1908 135
rect 1903 128 1905 130
rect 1907 128 1908 130
rect 1903 126 1908 128
rect 1903 119 1907 126
rect 1903 117 1904 119
rect 1906 117 1907 119
rect 1903 106 1907 117
rect 1935 131 1939 138
rect 1944 131 1949 140
rect 1935 129 1949 131
rect 1926 128 1949 129
rect 1926 126 1932 128
rect 1934 126 1946 128
rect 1948 126 1949 128
rect 1926 125 1939 126
rect 1943 125 1949 126
rect 1944 124 1949 125
rect 1918 120 1932 121
rect 1918 118 1922 120
rect 1924 118 1932 120
rect 1918 117 1932 118
rect 1903 104 1905 106
rect 1907 104 1915 106
rect 1903 100 1915 104
rect 1927 111 1932 117
rect 1927 109 1928 111
rect 1930 109 1932 111
rect 1927 108 1932 109
rect 1960 115 1965 122
rect 1988 137 2004 138
rect 1988 135 1990 137
rect 1992 135 2004 137
rect 1988 133 2004 135
rect 1960 114 1962 115
rect 1952 113 1962 114
rect 1964 113 1965 115
rect 1952 111 1965 113
rect 1952 109 1955 111
rect 1957 109 1965 111
rect 1952 108 1965 109
rect 2000 108 2004 133
rect 2000 106 2001 108
rect 2003 106 2004 108
rect 2000 105 2004 106
rect 1980 104 2004 105
rect 1980 102 1982 104
rect 1984 102 2004 104
rect 1980 101 2004 102
rect 771 94 2008 95
rect 23 92 36 94
rect 38 92 46 94
rect 48 92 94 94
rect 96 92 104 94
rect 106 92 116 94
rect 118 92 126 94
rect 128 92 157 94
rect 159 92 210 94
rect 212 92 240 94
rect 242 92 250 94
rect 252 92 281 94
rect 283 92 334 94
rect 336 93 778 94
rect 336 92 384 93
rect 23 91 384 92
rect 386 91 394 93
rect 396 91 424 93
rect 426 91 434 93
rect 436 91 452 93
rect 454 91 505 93
rect 507 91 536 93
rect 538 91 546 93
rect 548 91 589 93
rect 591 91 599 93
rect 601 91 629 93
rect 631 91 639 93
rect 641 91 657 93
rect 659 91 710 93
rect 712 91 741 93
rect 743 91 751 93
rect 753 92 778 93
rect 780 92 818 94
rect 820 92 828 94
rect 830 92 859 94
rect 861 92 912 94
rect 914 92 923 94
rect 925 92 933 94
rect 935 92 964 94
rect 966 92 1017 94
rect 1019 92 1028 94
rect 1030 92 1068 94
rect 1070 92 1078 94
rect 1080 92 1109 94
rect 1111 92 1162 94
rect 1164 92 1173 94
rect 1175 92 1183 94
rect 1185 92 1214 94
rect 1216 92 1267 94
rect 1269 92 1278 94
rect 1280 92 1318 94
rect 1320 92 1328 94
rect 1330 92 1359 94
rect 1361 92 1412 94
rect 1414 92 1423 94
rect 1425 92 1433 94
rect 1435 92 1464 94
rect 1466 92 1517 94
rect 1519 92 1528 94
rect 1530 92 1568 94
rect 1570 92 1578 94
rect 1580 92 1609 94
rect 1611 92 1662 94
rect 1664 92 1673 94
rect 1675 92 1683 94
rect 1685 92 1714 94
rect 1716 92 1767 94
rect 1769 92 1826 94
rect 1828 92 1836 94
rect 1838 92 1884 94
rect 1886 92 1894 94
rect 1896 92 1906 94
rect 1908 92 1916 94
rect 1918 92 1947 94
rect 1949 92 2000 94
rect 2002 92 2008 94
rect 753 91 2008 92
rect 23 88 2008 91
rect 23 87 756 88
rect 771 87 1775 88
rect 1813 87 2008 88
rect 353 86 756 87
rect 1031 86 1431 87
rect 436 77 441 86
rect 3 73 2017 77
rect 3 72 939 73
rect 3 70 10 72
rect 12 70 50 72
rect 52 70 60 72
rect 62 70 91 72
rect 93 70 144 72
rect 146 70 155 72
rect 157 70 165 72
rect 167 70 196 72
rect 198 70 249 72
rect 251 70 260 72
rect 262 70 300 72
rect 302 70 310 72
rect 312 70 341 72
rect 343 70 394 72
rect 396 70 405 72
rect 407 70 415 72
rect 417 70 446 72
rect 448 70 499 72
rect 501 70 510 72
rect 512 70 550 72
rect 552 70 560 72
rect 562 70 591 72
rect 593 70 644 72
rect 646 70 655 72
rect 657 70 665 72
rect 667 70 696 72
rect 698 70 749 72
rect 751 70 760 72
rect 762 70 800 72
rect 802 70 810 72
rect 812 70 841 72
rect 843 70 894 72
rect 896 70 905 72
rect 907 70 915 72
rect 917 71 939 72
rect 941 72 1110 73
rect 941 71 946 72
rect 917 70 946 71
rect 948 70 999 72
rect 1001 70 1020 72
rect 1022 70 1060 72
rect 1062 70 1070 72
rect 1072 70 1101 72
rect 1103 71 1110 72
rect 1112 72 1949 73
rect 1112 71 1154 72
rect 1103 70 1154 71
rect 1156 70 1165 72
rect 1167 70 1175 72
rect 1177 70 1206 72
rect 1208 70 1259 72
rect 1261 70 1270 72
rect 1272 70 1310 72
rect 1312 70 1320 72
rect 1322 70 1351 72
rect 1353 70 1360 72
rect 1362 70 1404 72
rect 1406 70 1415 72
rect 1417 70 1425 72
rect 1427 70 1456 72
rect 1458 70 1509 72
rect 1511 70 1520 72
rect 1522 70 1560 72
rect 1562 70 1570 72
rect 1572 70 1601 72
rect 1603 70 1654 72
rect 1656 70 1665 72
rect 1667 70 1675 72
rect 1677 70 1706 72
rect 1708 70 1759 72
rect 1761 70 1770 72
rect 1772 70 1810 72
rect 1812 70 1820 72
rect 1822 70 1851 72
rect 1853 70 1904 72
rect 1906 70 1915 72
rect 1917 70 1925 72
rect 1927 71 1949 72
rect 1951 72 2017 73
rect 1951 71 1956 72
rect 1927 70 1956 71
rect 1958 70 2009 72
rect 2011 70 2017 72
rect 3 69 2017 70
rect 47 60 59 64
rect 47 58 49 60
rect 51 58 59 60
rect 124 62 148 63
rect 7 55 12 57
rect 7 53 9 55
rect 11 53 12 55
rect 7 51 12 53
rect 7 32 11 51
rect 39 47 43 56
rect 47 47 51 58
rect 124 60 126 62
rect 128 60 148 62
rect 124 59 148 60
rect 7 30 9 32
rect 7 25 11 30
rect 7 23 9 25
rect 22 46 51 47
rect 22 44 26 46
rect 28 44 51 46
rect 22 43 51 44
rect 22 37 36 39
rect 38 37 43 39
rect 22 35 43 37
rect 39 29 43 35
rect 39 27 40 29
rect 42 27 43 29
rect 39 26 43 27
rect 47 38 51 43
rect 71 55 76 56
rect 71 53 72 55
rect 74 53 76 55
rect 71 47 76 53
rect 47 36 52 38
rect 47 34 49 36
rect 51 34 52 36
rect 47 29 52 34
rect 47 27 49 29
rect 51 27 52 29
rect 62 46 76 47
rect 62 44 66 46
rect 68 44 76 46
rect 62 43 76 44
rect 96 55 109 56
rect 96 53 99 55
rect 101 53 109 55
rect 96 51 109 53
rect 144 55 148 59
rect 96 50 106 51
rect 104 49 106 50
rect 108 49 109 51
rect 88 39 93 40
rect 70 38 83 39
rect 87 38 93 39
rect 70 36 71 38
rect 73 36 76 38
rect 78 36 90 38
rect 92 36 93 38
rect 70 35 93 36
rect 79 33 93 35
rect 104 42 109 49
rect 144 53 145 55
rect 147 53 148 55
rect 47 25 52 27
rect 7 19 20 23
rect 7 18 11 19
rect 79 26 83 33
rect 88 24 93 33
rect 88 18 100 24
rect 144 31 148 53
rect 132 29 148 31
rect 132 27 134 29
rect 136 27 148 29
rect 132 26 148 27
rect 152 60 164 64
rect 152 58 154 60
rect 156 58 164 60
rect 229 62 253 63
rect 152 38 156 58
rect 229 60 231 62
rect 233 60 253 62
rect 229 59 253 60
rect 176 55 181 56
rect 176 53 177 55
rect 179 53 181 55
rect 176 47 181 53
rect 152 36 157 38
rect 152 34 154 36
rect 156 34 157 36
rect 152 29 157 34
rect 152 27 154 29
rect 156 27 157 29
rect 167 46 181 47
rect 167 44 171 46
rect 173 44 181 46
rect 167 43 181 44
rect 201 55 214 56
rect 201 53 204 55
rect 206 53 214 55
rect 201 51 214 53
rect 201 50 211 51
rect 209 49 211 50
rect 213 49 214 51
rect 193 39 198 40
rect 175 38 188 39
rect 192 38 198 39
rect 175 36 181 38
rect 183 37 195 38
rect 183 36 187 37
rect 175 35 187 36
rect 189 36 195 37
rect 197 36 198 38
rect 189 35 198 36
rect 184 33 198 35
rect 209 42 214 49
rect 152 25 157 27
rect 184 26 188 33
rect 193 24 198 33
rect 193 18 205 24
rect 249 31 253 59
rect 297 60 309 64
rect 297 58 299 60
rect 301 58 309 60
rect 374 62 398 63
rect 237 29 253 31
rect 237 27 239 29
rect 241 27 253 29
rect 237 26 253 27
rect 257 55 262 57
rect 257 53 259 55
rect 261 53 262 55
rect 257 51 262 53
rect 257 37 261 51
rect 257 35 258 37
rect 260 35 261 37
rect 257 32 261 35
rect 289 47 293 56
rect 297 47 301 58
rect 374 60 376 62
rect 378 60 398 62
rect 374 59 398 60
rect 257 30 259 32
rect 257 25 261 30
rect 257 23 259 25
rect 272 46 301 47
rect 272 44 276 46
rect 278 44 301 46
rect 272 43 301 44
rect 272 37 286 39
rect 288 37 293 39
rect 272 35 293 37
rect 289 29 293 35
rect 289 27 290 29
rect 292 27 293 29
rect 289 26 293 27
rect 297 38 301 43
rect 321 55 326 56
rect 321 53 322 55
rect 324 53 326 55
rect 321 47 326 53
rect 297 36 302 38
rect 297 34 299 36
rect 301 34 302 36
rect 297 29 302 34
rect 297 27 299 29
rect 301 27 302 29
rect 312 46 326 47
rect 312 44 316 46
rect 318 44 326 46
rect 312 43 326 44
rect 346 55 359 56
rect 346 53 349 55
rect 351 53 359 55
rect 346 51 359 53
rect 394 55 398 59
rect 346 50 356 51
rect 354 49 356 50
rect 358 49 359 51
rect 338 39 343 40
rect 320 38 333 39
rect 337 38 343 39
rect 320 36 321 38
rect 323 36 326 38
rect 328 36 340 38
rect 342 36 343 38
rect 320 35 343 36
rect 329 33 343 35
rect 354 42 359 49
rect 394 53 395 55
rect 397 53 398 55
rect 297 25 302 27
rect 257 19 270 23
rect 257 18 261 19
rect 329 26 333 33
rect 338 24 343 33
rect 338 18 350 24
rect 394 31 398 53
rect 382 29 398 31
rect 382 27 384 29
rect 386 27 398 29
rect 382 26 398 27
rect 402 60 414 64
rect 402 58 404 60
rect 406 58 414 60
rect 479 62 503 63
rect 402 38 406 58
rect 479 60 481 62
rect 483 60 503 62
rect 479 59 503 60
rect 426 55 431 56
rect 426 53 427 55
rect 429 53 431 55
rect 426 47 431 53
rect 402 36 407 38
rect 402 34 404 36
rect 406 34 407 36
rect 402 29 407 34
rect 402 27 404 29
rect 406 27 407 29
rect 417 46 431 47
rect 417 44 421 46
rect 423 44 431 46
rect 417 43 431 44
rect 451 55 464 56
rect 451 53 454 55
rect 456 53 464 55
rect 451 51 464 53
rect 451 50 461 51
rect 459 49 461 50
rect 463 49 464 51
rect 443 39 448 40
rect 425 38 438 39
rect 442 38 448 39
rect 425 36 431 38
rect 433 37 445 38
rect 433 36 439 37
rect 425 35 439 36
rect 441 36 445 37
rect 447 36 448 38
rect 441 35 448 36
rect 434 33 448 35
rect 459 42 464 49
rect 402 25 407 27
rect 434 26 438 33
rect 443 24 448 33
rect 443 18 455 24
rect 499 31 503 59
rect 547 60 559 64
rect 547 58 549 60
rect 551 58 559 60
rect 624 62 648 63
rect 487 29 503 31
rect 487 27 489 29
rect 491 27 503 29
rect 487 26 503 27
rect 507 55 512 57
rect 507 53 509 55
rect 511 53 512 55
rect 507 51 512 53
rect 507 37 511 51
rect 507 35 508 37
rect 510 35 511 37
rect 507 32 511 35
rect 539 47 543 56
rect 547 47 551 58
rect 624 60 626 62
rect 628 60 648 62
rect 624 59 648 60
rect 507 30 509 32
rect 507 25 511 30
rect 507 23 509 25
rect 522 46 551 47
rect 522 44 526 46
rect 528 44 551 46
rect 522 43 551 44
rect 522 37 536 39
rect 538 37 543 39
rect 522 35 543 37
rect 539 29 543 35
rect 539 27 540 29
rect 542 27 543 29
rect 539 26 543 27
rect 547 38 551 43
rect 571 55 576 56
rect 571 53 572 55
rect 574 53 576 55
rect 571 47 576 53
rect 547 36 552 38
rect 547 34 549 36
rect 551 34 552 36
rect 547 29 552 34
rect 547 27 549 29
rect 551 27 552 29
rect 562 46 576 47
rect 562 44 566 46
rect 568 44 576 46
rect 562 43 576 44
rect 596 55 609 56
rect 596 53 599 55
rect 601 53 609 55
rect 596 51 609 53
rect 644 55 648 59
rect 596 50 606 51
rect 604 49 606 50
rect 608 49 609 51
rect 588 39 593 40
rect 570 38 583 39
rect 587 38 593 39
rect 570 36 576 38
rect 578 36 590 38
rect 592 36 593 38
rect 570 35 593 36
rect 579 33 593 35
rect 604 42 609 49
rect 644 53 645 55
rect 647 53 648 55
rect 547 25 552 27
rect 507 19 520 23
rect 507 18 511 19
rect 579 26 583 33
rect 588 24 593 33
rect 588 21 600 24
rect 588 19 597 21
rect 599 19 600 21
rect 588 18 600 19
rect 644 31 648 53
rect 632 29 648 31
rect 632 27 634 29
rect 636 27 648 29
rect 632 26 648 27
rect 652 60 664 64
rect 652 58 654 60
rect 656 58 664 60
rect 729 62 753 63
rect 652 38 656 58
rect 729 60 731 62
rect 733 60 753 62
rect 729 59 753 60
rect 676 55 681 56
rect 676 53 677 55
rect 679 53 681 55
rect 676 47 681 53
rect 652 36 657 38
rect 652 34 654 36
rect 656 34 657 36
rect 652 29 657 34
rect 652 27 654 29
rect 656 27 657 29
rect 667 46 681 47
rect 667 44 671 46
rect 673 44 681 46
rect 667 43 681 44
rect 701 55 714 56
rect 701 53 704 55
rect 706 53 714 55
rect 701 51 714 53
rect 701 50 711 51
rect 709 49 711 50
rect 713 49 714 51
rect 693 39 698 40
rect 675 38 688 39
rect 692 38 698 39
rect 675 36 681 38
rect 683 37 695 38
rect 683 36 689 37
rect 675 35 689 36
rect 691 36 695 37
rect 697 36 698 38
rect 691 35 698 36
rect 684 33 698 35
rect 709 42 714 49
rect 652 25 657 27
rect 684 26 688 33
rect 693 24 698 33
rect 693 18 705 24
rect 749 31 753 59
rect 797 60 809 64
rect 797 58 799 60
rect 801 58 809 60
rect 874 62 898 63
rect 737 29 753 31
rect 737 27 739 29
rect 741 27 753 29
rect 737 26 753 27
rect 757 55 762 57
rect 757 53 759 55
rect 761 53 762 55
rect 757 51 762 53
rect 757 37 761 51
rect 757 35 758 37
rect 760 35 761 37
rect 757 32 761 35
rect 789 47 793 56
rect 797 47 801 58
rect 874 60 876 62
rect 878 60 898 62
rect 874 59 898 60
rect 757 30 759 32
rect 757 25 761 30
rect 757 23 759 25
rect 772 46 801 47
rect 772 44 776 46
rect 778 44 801 46
rect 772 43 801 44
rect 772 37 786 39
rect 788 37 793 39
rect 772 35 793 37
rect 789 29 793 35
rect 789 27 790 29
rect 792 27 793 29
rect 789 26 793 27
rect 797 38 801 43
rect 821 55 826 56
rect 821 53 822 55
rect 824 53 826 55
rect 821 47 826 53
rect 797 36 802 38
rect 797 34 799 36
rect 801 34 802 36
rect 797 29 802 34
rect 797 27 799 29
rect 801 27 802 29
rect 812 46 826 47
rect 812 44 816 46
rect 818 44 826 46
rect 812 43 826 44
rect 846 55 859 56
rect 846 53 849 55
rect 851 53 859 55
rect 846 51 859 53
rect 894 55 898 59
rect 846 50 856 51
rect 854 49 856 50
rect 858 49 859 51
rect 838 39 843 40
rect 820 38 833 39
rect 837 38 843 39
rect 820 36 826 38
rect 828 36 840 38
rect 842 36 843 38
rect 820 35 843 36
rect 829 33 843 35
rect 854 45 859 49
rect 894 53 895 55
rect 897 53 898 55
rect 854 43 856 45
rect 858 43 859 45
rect 854 42 859 43
rect 797 25 802 27
rect 757 19 770 23
rect 757 18 761 19
rect 829 26 833 33
rect 838 24 843 33
rect 838 21 850 24
rect 838 19 847 21
rect 849 19 850 21
rect 838 18 850 19
rect 894 31 898 53
rect 882 29 898 31
rect 882 27 884 29
rect 886 27 898 29
rect 882 26 898 27
rect 902 60 914 64
rect 902 58 904 60
rect 906 58 914 60
rect 979 62 1003 63
rect 902 38 906 58
rect 979 60 981 62
rect 983 60 1003 62
rect 979 59 1003 60
rect 926 55 931 56
rect 926 53 927 55
rect 929 53 931 55
rect 926 47 931 53
rect 902 36 907 38
rect 902 34 904 36
rect 906 34 907 36
rect 902 29 907 34
rect 902 27 904 29
rect 906 27 907 29
rect 917 46 931 47
rect 917 44 921 46
rect 923 44 931 46
rect 917 43 931 44
rect 951 55 964 56
rect 951 53 954 55
rect 956 53 964 55
rect 951 51 964 53
rect 951 50 961 51
rect 959 49 961 50
rect 963 49 964 51
rect 943 39 948 40
rect 925 38 948 39
rect 925 36 931 38
rect 933 36 939 38
rect 941 36 945 38
rect 947 36 948 38
rect 925 35 948 36
rect 934 33 948 35
rect 959 42 964 49
rect 902 25 907 27
rect 934 26 938 33
rect 943 24 948 33
rect 943 18 955 24
rect 999 31 1003 59
rect 1057 60 1069 64
rect 1057 58 1059 60
rect 1061 58 1069 60
rect 1134 62 1158 63
rect 987 29 1003 31
rect 987 27 989 29
rect 991 27 1003 29
rect 987 26 1003 27
rect 1017 55 1022 57
rect 1017 53 1019 55
rect 1021 53 1022 55
rect 1017 51 1022 53
rect 1017 32 1021 51
rect 1049 47 1053 56
rect 1057 47 1061 58
rect 1134 60 1136 62
rect 1138 60 1158 62
rect 1134 59 1158 60
rect 1017 30 1019 32
rect 1017 25 1021 30
rect 1017 23 1019 25
rect 1032 46 1061 47
rect 1032 44 1036 46
rect 1038 44 1061 46
rect 1032 43 1061 44
rect 1032 37 1046 39
rect 1048 37 1053 39
rect 1032 35 1053 37
rect 1049 29 1053 35
rect 1049 27 1050 29
rect 1052 27 1053 29
rect 1049 26 1053 27
rect 1057 38 1061 43
rect 1081 55 1086 56
rect 1081 53 1082 55
rect 1084 53 1086 55
rect 1081 47 1086 53
rect 1057 36 1062 38
rect 1057 34 1059 36
rect 1061 34 1062 36
rect 1057 29 1062 34
rect 1057 27 1059 29
rect 1061 27 1062 29
rect 1072 46 1086 47
rect 1072 44 1076 46
rect 1078 44 1086 46
rect 1072 43 1086 44
rect 1106 55 1119 56
rect 1106 53 1109 55
rect 1111 53 1119 55
rect 1106 51 1119 53
rect 1154 55 1158 59
rect 1106 50 1116 51
rect 1114 49 1116 50
rect 1118 49 1119 51
rect 1098 39 1103 40
rect 1080 38 1093 39
rect 1097 38 1103 39
rect 1080 36 1086 38
rect 1088 37 1100 38
rect 1088 36 1094 37
rect 1080 35 1094 36
rect 1096 36 1100 37
rect 1102 36 1103 38
rect 1096 35 1103 36
rect 1089 33 1103 35
rect 1114 42 1119 49
rect 1154 53 1155 55
rect 1157 53 1158 55
rect 1057 25 1062 27
rect 1017 19 1030 23
rect 1017 18 1021 19
rect 1089 26 1093 33
rect 1098 24 1103 33
rect 1098 18 1110 24
rect 1154 31 1158 53
rect 1142 29 1158 31
rect 1142 27 1144 29
rect 1146 27 1158 29
rect 1142 26 1158 27
rect 1162 60 1174 64
rect 1162 58 1164 60
rect 1166 58 1174 60
rect 1239 62 1263 63
rect 1162 38 1166 58
rect 1239 60 1241 62
rect 1243 60 1245 62
rect 1247 60 1263 62
rect 1239 59 1263 60
rect 1186 55 1191 56
rect 1186 53 1187 55
rect 1189 53 1191 55
rect 1186 47 1191 53
rect 1162 36 1167 38
rect 1162 34 1164 36
rect 1166 34 1167 36
rect 1162 29 1167 34
rect 1162 27 1164 29
rect 1166 27 1167 29
rect 1177 46 1191 47
rect 1177 44 1181 46
rect 1183 44 1191 46
rect 1177 43 1191 44
rect 1211 55 1224 56
rect 1211 53 1214 55
rect 1216 53 1224 55
rect 1211 51 1224 53
rect 1211 50 1221 51
rect 1219 49 1221 50
rect 1223 49 1224 51
rect 1203 39 1208 40
rect 1185 38 1198 39
rect 1202 38 1208 39
rect 1185 36 1191 38
rect 1193 37 1205 38
rect 1193 36 1197 37
rect 1185 35 1197 36
rect 1199 36 1205 37
rect 1207 36 1208 38
rect 1199 35 1208 36
rect 1194 33 1208 35
rect 1219 42 1224 49
rect 1162 25 1167 27
rect 1194 26 1198 33
rect 1203 24 1208 33
rect 1203 18 1215 24
rect 1259 31 1263 59
rect 1307 60 1319 64
rect 1307 58 1309 60
rect 1311 58 1319 60
rect 1384 62 1408 63
rect 1247 29 1263 31
rect 1247 27 1249 29
rect 1251 27 1263 29
rect 1247 26 1263 27
rect 1267 55 1272 57
rect 1267 53 1269 55
rect 1271 53 1272 55
rect 1267 51 1272 53
rect 1267 37 1271 51
rect 1267 35 1268 37
rect 1270 35 1271 37
rect 1267 32 1271 35
rect 1299 47 1303 56
rect 1307 47 1311 58
rect 1384 60 1386 62
rect 1388 60 1408 62
rect 1384 59 1408 60
rect 1267 30 1269 32
rect 1267 25 1271 30
rect 1267 23 1269 25
rect 1282 46 1311 47
rect 1282 44 1286 46
rect 1288 44 1311 46
rect 1282 43 1311 44
rect 1282 37 1296 39
rect 1298 37 1303 39
rect 1282 35 1303 37
rect 1299 29 1303 35
rect 1299 27 1300 29
rect 1302 27 1303 29
rect 1299 26 1303 27
rect 1307 38 1311 43
rect 1331 55 1336 56
rect 1331 53 1332 55
rect 1334 53 1336 55
rect 1331 47 1336 53
rect 1307 36 1312 38
rect 1307 34 1309 36
rect 1311 34 1312 36
rect 1307 29 1312 34
rect 1307 27 1309 29
rect 1311 27 1312 29
rect 1322 46 1336 47
rect 1322 44 1326 46
rect 1328 44 1336 46
rect 1322 43 1336 44
rect 1356 55 1369 56
rect 1356 53 1359 55
rect 1361 53 1369 55
rect 1356 51 1369 53
rect 1404 55 1408 59
rect 1356 50 1366 51
rect 1364 49 1366 50
rect 1368 49 1369 51
rect 1348 39 1353 40
rect 1330 38 1353 39
rect 1330 36 1336 38
rect 1338 37 1350 38
rect 1338 36 1345 37
rect 1330 35 1345 36
rect 1347 36 1350 37
rect 1352 36 1353 38
rect 1347 35 1353 36
rect 1339 33 1353 35
rect 1364 42 1369 49
rect 1404 53 1405 55
rect 1407 53 1408 55
rect 1307 25 1312 27
rect 1267 19 1280 23
rect 1267 18 1271 19
rect 1339 26 1343 33
rect 1348 24 1353 33
rect 1348 18 1360 24
rect 1404 31 1408 53
rect 1392 29 1408 31
rect 1392 27 1394 29
rect 1396 27 1408 29
rect 1392 26 1408 27
rect 1412 60 1424 64
rect 1412 58 1414 60
rect 1416 58 1424 60
rect 1489 62 1513 63
rect 1412 38 1416 58
rect 1489 60 1491 62
rect 1493 60 1513 62
rect 1489 59 1513 60
rect 1436 55 1441 56
rect 1436 53 1437 55
rect 1439 53 1441 55
rect 1436 47 1441 53
rect 1412 36 1417 38
rect 1412 34 1414 36
rect 1416 34 1417 36
rect 1412 29 1417 34
rect 1412 27 1414 29
rect 1416 27 1417 29
rect 1427 46 1441 47
rect 1427 44 1431 46
rect 1433 44 1441 46
rect 1427 43 1441 44
rect 1461 55 1474 56
rect 1461 53 1464 55
rect 1466 53 1474 55
rect 1461 51 1474 53
rect 1461 50 1471 51
rect 1469 49 1471 50
rect 1473 49 1474 51
rect 1453 39 1458 40
rect 1435 38 1448 39
rect 1452 38 1458 39
rect 1435 36 1441 38
rect 1443 37 1455 38
rect 1443 36 1449 37
rect 1435 35 1449 36
rect 1451 36 1455 37
rect 1457 36 1458 38
rect 1451 35 1458 36
rect 1444 33 1458 35
rect 1469 42 1474 49
rect 1509 45 1513 59
rect 1557 60 1569 64
rect 1557 58 1559 60
rect 1561 58 1569 60
rect 1634 62 1658 63
rect 1509 43 1510 45
rect 1512 43 1513 45
rect 1412 25 1417 27
rect 1444 26 1448 33
rect 1453 24 1458 33
rect 1453 18 1465 24
rect 1509 31 1513 43
rect 1497 29 1513 31
rect 1497 27 1499 29
rect 1501 27 1513 29
rect 1497 26 1513 27
rect 1517 55 1522 57
rect 1517 53 1519 55
rect 1521 53 1522 55
rect 1517 51 1522 53
rect 1517 37 1521 51
rect 1517 35 1518 37
rect 1520 35 1521 37
rect 1517 32 1521 35
rect 1549 47 1553 56
rect 1557 47 1561 58
rect 1634 60 1636 62
rect 1638 60 1658 62
rect 1634 59 1658 60
rect 1517 30 1519 32
rect 1517 25 1521 30
rect 1517 23 1519 25
rect 1532 46 1561 47
rect 1532 44 1536 46
rect 1538 44 1561 46
rect 1532 43 1561 44
rect 1532 37 1546 39
rect 1548 37 1553 39
rect 1532 35 1553 37
rect 1549 29 1553 35
rect 1549 27 1550 29
rect 1552 27 1553 29
rect 1549 26 1553 27
rect 1557 38 1561 43
rect 1581 55 1586 56
rect 1581 53 1582 55
rect 1584 53 1586 55
rect 1581 47 1586 53
rect 1557 36 1562 38
rect 1557 34 1559 36
rect 1561 34 1562 36
rect 1557 29 1562 34
rect 1557 27 1559 29
rect 1561 27 1562 29
rect 1572 46 1586 47
rect 1572 44 1576 46
rect 1578 44 1586 46
rect 1572 43 1586 44
rect 1606 55 1619 56
rect 1606 53 1609 55
rect 1611 53 1619 55
rect 1606 51 1619 53
rect 1654 55 1658 59
rect 1606 50 1616 51
rect 1614 49 1616 50
rect 1618 49 1619 51
rect 1598 39 1603 40
rect 1580 38 1603 39
rect 1580 36 1582 38
rect 1584 36 1586 38
rect 1588 36 1600 38
rect 1602 36 1603 38
rect 1580 35 1603 36
rect 1589 33 1603 35
rect 1614 42 1619 49
rect 1654 53 1655 55
rect 1657 53 1658 55
rect 1557 25 1562 27
rect 1517 19 1530 23
rect 1517 18 1521 19
rect 1589 26 1593 33
rect 1598 24 1603 33
rect 1598 18 1610 24
rect 1654 31 1658 53
rect 1642 29 1658 31
rect 1642 27 1644 29
rect 1646 27 1658 29
rect 1642 26 1658 27
rect 1662 60 1674 64
rect 1662 58 1664 60
rect 1666 58 1674 60
rect 1739 62 1763 63
rect 1662 38 1666 58
rect 1739 60 1741 62
rect 1743 60 1763 62
rect 1739 59 1763 60
rect 1686 55 1691 56
rect 1686 53 1687 55
rect 1689 53 1691 55
rect 1686 47 1691 53
rect 1662 36 1667 38
rect 1662 34 1664 36
rect 1666 34 1667 36
rect 1662 29 1667 34
rect 1662 27 1664 29
rect 1666 27 1667 29
rect 1677 46 1691 47
rect 1677 44 1681 46
rect 1683 44 1691 46
rect 1677 43 1691 44
rect 1711 55 1724 56
rect 1711 53 1714 55
rect 1716 53 1724 55
rect 1711 51 1724 53
rect 1711 50 1721 51
rect 1719 49 1721 50
rect 1723 49 1724 51
rect 1703 39 1708 40
rect 1685 38 1698 39
rect 1702 38 1708 39
rect 1685 36 1691 38
rect 1693 37 1705 38
rect 1693 36 1699 37
rect 1685 35 1699 36
rect 1701 36 1705 37
rect 1707 36 1708 38
rect 1701 35 1708 36
rect 1694 33 1708 35
rect 1719 42 1724 49
rect 1662 25 1667 27
rect 1694 26 1698 33
rect 1703 24 1708 33
rect 1703 18 1715 24
rect 1759 31 1763 59
rect 1807 60 1819 64
rect 1807 58 1809 60
rect 1811 58 1819 60
rect 1884 62 1908 63
rect 1747 29 1763 31
rect 1747 27 1749 29
rect 1751 27 1763 29
rect 1747 26 1763 27
rect 1767 55 1772 57
rect 1767 53 1769 55
rect 1771 53 1772 55
rect 1767 51 1772 53
rect 1767 37 1771 51
rect 1767 35 1768 37
rect 1770 35 1771 37
rect 1767 32 1771 35
rect 1799 47 1803 56
rect 1807 47 1811 58
rect 1884 60 1886 62
rect 1888 60 1908 62
rect 1884 59 1908 60
rect 1767 30 1769 32
rect 1767 25 1771 30
rect 1767 23 1769 25
rect 1782 46 1811 47
rect 1782 44 1786 46
rect 1788 44 1811 46
rect 1782 43 1811 44
rect 1782 37 1796 39
rect 1798 37 1803 39
rect 1782 35 1803 37
rect 1799 29 1803 35
rect 1799 27 1800 29
rect 1802 27 1803 29
rect 1799 26 1803 27
rect 1807 38 1811 43
rect 1831 55 1836 56
rect 1831 53 1832 55
rect 1834 53 1836 55
rect 1831 47 1836 53
rect 1807 36 1812 38
rect 1807 34 1809 36
rect 1811 34 1812 36
rect 1807 29 1812 34
rect 1807 27 1809 29
rect 1811 27 1812 29
rect 1822 46 1836 47
rect 1822 44 1826 46
rect 1828 44 1836 46
rect 1822 43 1836 44
rect 1856 55 1869 56
rect 1856 53 1859 55
rect 1861 53 1869 55
rect 1856 51 1869 53
rect 1904 55 1908 59
rect 1856 50 1866 51
rect 1864 49 1866 50
rect 1868 49 1869 51
rect 1848 39 1853 40
rect 1830 38 1853 39
rect 1830 36 1832 38
rect 1834 36 1836 38
rect 1838 36 1850 38
rect 1852 36 1853 38
rect 1830 35 1853 36
rect 1839 33 1853 35
rect 1864 42 1869 49
rect 1904 53 1905 55
rect 1907 53 1908 55
rect 1807 25 1812 27
rect 1767 19 1780 23
rect 1767 18 1771 19
rect 1839 26 1843 33
rect 1848 24 1853 33
rect 1848 18 1860 24
rect 1904 31 1908 53
rect 1892 29 1908 31
rect 1892 27 1894 29
rect 1896 27 1908 29
rect 1892 26 1908 27
rect 1912 60 1924 64
rect 1912 58 1914 60
rect 1916 58 1924 60
rect 1989 62 2013 63
rect 1912 38 1916 58
rect 1989 60 1991 62
rect 1993 60 2013 62
rect 1989 59 2013 60
rect 1936 55 1941 56
rect 1936 53 1937 55
rect 1939 53 1941 55
rect 1936 47 1941 53
rect 1912 36 1917 38
rect 1912 34 1914 36
rect 1916 34 1917 36
rect 1912 29 1917 34
rect 1912 27 1914 29
rect 1916 27 1917 29
rect 1927 46 1941 47
rect 1927 44 1931 46
rect 1933 44 1941 46
rect 1927 43 1941 44
rect 1961 55 1974 56
rect 1961 53 1964 55
rect 1966 53 1974 55
rect 1961 51 1974 53
rect 1961 50 1971 51
rect 1969 49 1971 50
rect 1973 49 1974 51
rect 1953 39 1958 40
rect 1935 38 1958 39
rect 1935 36 1941 38
rect 1943 36 1949 38
rect 1951 36 1955 38
rect 1957 36 1958 38
rect 1935 35 1958 36
rect 1944 33 1958 35
rect 1969 42 1974 49
rect 1912 25 1917 27
rect 1944 26 1948 33
rect 1953 24 1958 33
rect 1953 18 1965 24
rect 2009 31 2013 59
rect 1997 29 2013 31
rect 1997 27 1999 29
rect 2001 27 2013 29
rect 1997 26 2013 27
rect 3 12 2017 13
rect 3 10 10 12
rect 12 10 50 12
rect 52 10 124 12
rect 126 10 155 12
rect 157 10 229 12
rect 231 10 260 12
rect 262 10 300 12
rect 302 10 374 12
rect 376 10 405 12
rect 407 10 479 12
rect 481 10 510 12
rect 512 10 550 12
rect 552 10 624 12
rect 626 10 655 12
rect 657 10 729 12
rect 731 10 760 12
rect 762 10 800 12
rect 802 10 874 12
rect 876 10 905 12
rect 907 10 979 12
rect 981 10 1020 12
rect 1022 10 1060 12
rect 1062 10 1134 12
rect 1136 10 1165 12
rect 1167 10 1239 12
rect 1241 10 1270 12
rect 1272 10 1310 12
rect 1312 10 1384 12
rect 1386 10 1415 12
rect 1417 10 1489 12
rect 1491 10 1520 12
rect 1522 10 1560 12
rect 1562 10 1634 12
rect 1636 10 1665 12
rect 1667 10 1739 12
rect 1741 10 1770 12
rect 1772 10 1810 12
rect 1812 10 1884 12
rect 1886 10 1915 12
rect 1917 10 1989 12
rect 1991 10 2017 12
rect 3 5 2017 10
<< alu2 >>
rect 443 225 868 230
rect 443 221 448 225
rect 443 219 445 221
rect 447 219 448 221
rect 443 214 448 219
rect 355 210 407 214
rect 540 212 544 221
rect 560 210 612 214
rect 65 209 197 210
rect 65 207 66 209
rect 68 207 167 209
rect 169 207 194 209
rect 196 207 197 209
rect 65 206 197 207
rect 48 200 54 201
rect 48 198 51 200
rect 53 198 54 200
rect 25 184 37 185
rect 25 182 34 184
rect 36 182 37 184
rect 25 180 37 182
rect 25 107 30 180
rect 34 121 38 122
rect 34 119 35 121
rect 37 119 38 121
rect 34 116 38 119
rect 48 120 54 198
rect 90 200 94 201
rect 90 198 91 200
rect 93 198 94 200
rect 73 185 77 186
rect 73 183 74 185
rect 76 183 77 185
rect 73 159 77 183
rect 65 155 77 159
rect 65 137 69 155
rect 65 135 66 137
rect 68 135 69 137
rect 65 134 69 135
rect 48 118 49 120
rect 51 118 54 120
rect 48 117 54 118
rect 73 128 77 129
rect 73 126 74 128
rect 76 126 77 128
rect 34 114 35 116
rect 37 114 38 116
rect 34 113 38 114
rect 73 107 77 126
rect 90 120 94 198
rect 217 197 221 201
rect 120 194 124 197
rect 120 192 121 194
rect 123 192 124 194
rect 120 191 124 192
rect 217 195 218 197
rect 220 195 221 197
rect 104 186 189 187
rect 104 184 105 186
rect 107 184 186 186
rect 188 184 189 186
rect 104 183 189 184
rect 120 178 124 179
rect 120 176 121 178
rect 123 176 124 178
rect 120 160 124 176
rect 217 160 221 195
rect 120 159 130 160
rect 120 157 126 159
rect 128 157 130 159
rect 120 156 130 157
rect 161 155 221 160
rect 161 144 166 155
rect 161 142 162 144
rect 164 142 166 144
rect 161 140 166 142
rect 355 137 360 210
rect 364 204 368 206
rect 364 202 365 204
rect 367 202 368 204
rect 364 189 368 202
rect 364 187 365 189
rect 367 187 368 189
rect 364 186 368 187
rect 378 199 384 200
rect 378 197 379 199
rect 381 197 384 199
rect 355 135 367 137
rect 355 133 364 135
rect 366 133 367 135
rect 355 132 367 133
rect 90 118 91 120
rect 93 118 94 120
rect 90 117 94 118
rect 113 119 117 121
rect 113 117 114 119
rect 116 117 117 119
rect 113 116 117 117
rect 378 119 384 197
rect 403 191 407 210
rect 435 209 473 210
rect 435 208 500 209
rect 435 206 436 208
rect 438 206 468 208
rect 470 206 495 208
rect 497 206 500 208
rect 435 205 500 206
rect 443 200 448 201
rect 403 189 404 191
rect 406 189 407 191
rect 403 188 407 189
rect 420 199 424 200
rect 420 197 421 199
rect 423 197 424 199
rect 395 182 399 183
rect 395 180 396 182
rect 398 180 399 182
rect 395 162 399 180
rect 395 158 407 162
rect 403 134 407 158
rect 403 132 404 134
rect 406 132 407 134
rect 403 131 407 132
rect 378 117 381 119
rect 383 117 384 119
rect 378 116 384 117
rect 420 119 424 197
rect 443 198 444 200
rect 446 198 448 200
rect 443 193 448 198
rect 491 175 496 177
rect 491 173 492 175
rect 494 173 496 175
rect 491 162 496 173
rect 491 157 551 162
rect 434 133 519 134
rect 434 131 435 133
rect 437 131 516 133
rect 518 131 519 133
rect 434 130 519 131
rect 420 117 421 119
rect 423 117 424 119
rect 420 116 424 117
rect 547 122 551 157
rect 560 137 565 210
rect 583 199 589 200
rect 583 197 584 199
rect 586 197 589 199
rect 569 186 574 191
rect 569 184 570 186
rect 572 184 574 186
rect 569 178 574 184
rect 560 135 572 137
rect 560 133 569 135
rect 571 133 572 135
rect 560 132 572 133
rect 547 120 548 122
rect 550 120 551 122
rect 547 116 551 120
rect 583 119 589 197
rect 608 191 612 210
rect 640 209 678 210
rect 640 208 705 209
rect 640 206 641 208
rect 643 206 673 208
rect 675 206 700 208
rect 702 206 705 208
rect 640 205 705 206
rect 858 208 864 225
rect 858 206 860 208
rect 862 206 864 208
rect 1855 209 1987 210
rect 1855 207 1856 209
rect 1858 207 1957 209
rect 1959 207 1984 209
rect 1986 207 1987 209
rect 1855 206 1987 207
rect 858 204 864 206
rect 1838 200 1844 201
rect 608 189 609 191
rect 611 189 612 191
rect 608 188 612 189
rect 625 199 629 200
rect 625 197 626 199
rect 628 197 629 199
rect 600 182 604 183
rect 600 180 601 182
rect 603 180 604 182
rect 600 162 604 180
rect 600 158 612 162
rect 608 134 612 158
rect 608 132 609 134
rect 611 132 612 134
rect 608 131 612 132
rect 583 117 586 119
rect 588 117 589 119
rect 583 116 589 117
rect 625 119 629 197
rect 648 198 878 200
rect 648 196 649 198
rect 651 196 878 198
rect 648 195 875 196
rect 873 194 875 195
rect 877 194 878 196
rect 873 188 878 194
rect 1838 198 1841 200
rect 1843 198 1844 200
rect 1815 184 1827 185
rect 745 182 1041 184
rect 745 180 746 182
rect 748 180 1041 182
rect 745 179 1041 180
rect 696 175 701 177
rect 696 173 697 175
rect 699 173 701 175
rect 696 162 701 173
rect 873 170 878 173
rect 873 168 874 170
rect 876 168 878 170
rect 696 157 756 162
rect 639 133 724 134
rect 639 131 640 133
rect 642 131 721 133
rect 723 131 724 133
rect 639 130 724 131
rect 752 122 756 157
rect 873 147 878 168
rect 873 145 874 147
rect 876 145 878 147
rect 873 143 878 145
rect 807 137 925 138
rect 807 135 808 137
rect 810 135 922 137
rect 924 135 925 137
rect 807 134 925 135
rect 954 129 1029 130
rect 856 128 861 129
rect 856 126 858 128
rect 860 126 861 128
rect 954 127 955 129
rect 957 127 1026 129
rect 1028 127 1029 129
rect 954 126 1029 127
rect 856 124 861 126
rect 752 120 753 122
rect 755 120 756 122
rect 625 117 626 119
rect 628 117 629 119
rect 625 116 629 117
rect 655 118 659 119
rect 655 116 656 118
rect 658 116 659 118
rect 752 116 756 120
rect 873 123 878 125
rect 873 121 874 123
rect 876 121 878 123
rect 655 115 659 116
rect 873 112 878 121
rect 105 111 170 112
rect 105 109 106 111
rect 108 109 138 111
rect 140 109 165 111
rect 167 109 170 111
rect 105 108 170 109
rect 210 110 214 112
rect 210 108 211 110
rect 213 108 214 110
rect 105 107 143 108
rect 25 103 77 107
rect 210 92 214 108
rect 237 109 241 112
rect 237 107 238 109
rect 240 107 241 109
rect 261 111 294 112
rect 839 111 878 112
rect 261 109 262 111
rect 264 109 289 111
rect 291 109 294 111
rect 261 108 294 109
rect 395 110 527 111
rect 395 108 396 110
rect 398 108 497 110
rect 499 108 524 110
rect 526 108 527 110
rect 395 107 527 108
rect 600 110 732 111
rect 600 108 601 110
rect 603 108 702 110
rect 704 108 729 110
rect 731 108 732 110
rect 839 109 840 111
rect 842 109 867 111
rect 869 109 878 111
rect 839 108 878 109
rect 887 119 1028 121
rect 887 117 1018 119
rect 1020 117 1028 119
rect 887 116 1028 117
rect 600 107 732 108
rect 237 106 241 107
rect 29 91 40 92
rect 210 91 233 92
rect 29 89 35 91
rect 37 89 40 91
rect 29 88 40 89
rect 61 90 117 91
rect 61 88 114 90
rect 116 88 117 90
rect 210 89 221 91
rect 223 89 233 91
rect 210 88 233 89
rect 29 4 34 88
rect 61 87 117 88
rect 61 39 67 87
rect 237 82 242 106
rect 887 105 892 116
rect 1035 112 1041 179
rect 1815 182 1824 184
rect 1826 182 1827 184
rect 1815 180 1827 182
rect 1057 137 1175 138
rect 1057 135 1058 137
rect 1060 135 1172 137
rect 1174 135 1175 137
rect 1057 134 1175 135
rect 1307 137 1425 138
rect 1307 135 1308 137
rect 1310 135 1422 137
rect 1424 135 1425 137
rect 1307 134 1425 135
rect 1557 137 1675 138
rect 1557 135 1558 137
rect 1560 135 1672 137
rect 1674 135 1675 137
rect 1557 134 1675 135
rect 1206 129 1279 130
rect 1206 127 1207 129
rect 1209 127 1276 129
rect 1278 127 1279 129
rect 1206 126 1279 127
rect 1456 129 1529 130
rect 1456 127 1457 129
rect 1459 127 1526 129
rect 1528 127 1529 129
rect 1456 126 1529 127
rect 1606 128 1611 130
rect 1606 126 1608 128
rect 1610 126 1611 128
rect 1606 124 1611 126
rect 1045 119 1392 121
rect 1045 117 1049 119
rect 1051 117 1392 119
rect 1045 116 1392 117
rect 912 111 977 112
rect 912 109 913 111
rect 915 109 945 111
rect 947 109 972 111
rect 974 109 977 111
rect 1035 111 1122 112
rect 1035 110 1090 111
rect 912 108 977 109
rect 1036 109 1090 110
rect 1092 109 1117 111
rect 1119 109 1122 111
rect 1036 108 1122 109
rect 1162 111 1227 112
rect 1162 109 1163 111
rect 1165 109 1195 111
rect 1197 109 1222 111
rect 1224 109 1227 111
rect 1162 108 1227 109
rect 1339 111 1372 112
rect 1339 109 1340 111
rect 1342 109 1367 111
rect 1369 109 1372 111
rect 1339 108 1372 109
rect 334 104 338 105
rect 334 102 335 104
rect 337 102 338 104
rect 887 103 889 105
rect 891 103 892 105
rect 248 91 298 92
rect 248 89 256 91
rect 258 89 298 91
rect 248 88 298 89
rect 104 78 242 82
rect 104 56 108 78
rect 71 55 109 56
rect 71 53 72 55
rect 74 53 99 55
rect 101 53 109 55
rect 71 52 109 53
rect 144 55 209 56
rect 144 53 145 55
rect 147 53 177 55
rect 179 53 204 55
rect 206 53 209 55
rect 144 52 209 53
rect 294 39 298 88
rect 334 56 338 102
rect 655 101 659 102
rect 887 101 892 103
rect 1017 104 1021 106
rect 1017 102 1018 104
rect 1020 102 1021 104
rect 655 99 656 101
rect 658 99 659 101
rect 655 97 659 99
rect 655 95 1013 97
rect 655 93 1008 95
rect 1010 93 1013 95
rect 655 92 1013 93
rect 655 91 957 92
rect 1017 85 1021 102
rect 1267 105 1271 106
rect 1267 103 1268 105
rect 1270 103 1271 105
rect 1028 95 1101 97
rect 1028 93 1032 95
rect 1034 93 1101 95
rect 1028 92 1101 93
rect 1097 90 1263 92
rect 1097 88 1257 90
rect 1259 88 1263 90
rect 1097 87 1263 88
rect 928 79 956 83
rect 1017 80 1087 85
rect 1267 83 1271 103
rect 1339 92 1344 108
rect 1275 90 1344 92
rect 1275 88 1282 90
rect 1284 88 1344 90
rect 1386 95 1392 116
rect 1412 111 1477 112
rect 1412 109 1413 111
rect 1415 109 1445 111
rect 1447 109 1472 111
rect 1474 109 1477 111
rect 1412 108 1477 109
rect 1589 111 1622 112
rect 1589 109 1590 111
rect 1592 109 1617 111
rect 1619 109 1622 111
rect 1589 108 1622 109
rect 1662 111 1727 112
rect 1662 109 1663 111
rect 1665 109 1695 111
rect 1697 109 1722 111
rect 1724 109 1727 111
rect 1662 108 1727 109
rect 1517 105 1521 108
rect 1517 103 1518 105
rect 1520 103 1521 105
rect 1386 92 1510 95
rect 1386 90 1503 92
rect 1505 90 1510 92
rect 1386 89 1510 90
rect 1275 87 1344 88
rect 1517 85 1521 103
rect 1589 95 1594 108
rect 1815 107 1820 180
rect 1838 120 1844 198
rect 1880 200 1884 201
rect 1880 198 1881 200
rect 1883 198 1884 200
rect 1863 185 1867 186
rect 1863 183 1864 185
rect 1866 183 1867 185
rect 1863 159 1867 183
rect 1855 155 1867 159
rect 1855 137 1859 155
rect 1855 135 1856 137
rect 1858 135 1859 137
rect 1855 134 1859 135
rect 1838 118 1839 120
rect 1841 118 1844 120
rect 1838 117 1844 118
rect 1863 128 1867 129
rect 1863 126 1864 128
rect 1866 126 1867 128
rect 1863 107 1867 126
rect 1880 120 1884 198
rect 2007 197 2011 201
rect 2007 195 2008 197
rect 2010 195 2011 197
rect 1894 186 1979 187
rect 1894 184 1895 186
rect 1897 184 1976 186
rect 1978 184 1979 186
rect 1894 183 1979 184
rect 2007 160 2011 195
rect 1951 155 2011 160
rect 1951 144 1956 155
rect 1951 142 1952 144
rect 1954 142 1956 144
rect 1951 140 1956 142
rect 1880 118 1881 120
rect 1883 118 1884 120
rect 1880 117 1884 118
rect 1903 119 1907 120
rect 1903 117 1904 119
rect 1906 117 1907 119
rect 1903 116 1907 117
rect 1895 111 1960 112
rect 1895 109 1896 111
rect 1898 109 1928 111
rect 1930 109 1955 111
rect 1957 109 1960 111
rect 1895 108 1960 109
rect 2000 108 2004 110
rect 1895 107 1933 108
rect 1767 104 1804 105
rect 1767 102 1768 104
rect 1770 102 1804 104
rect 1815 103 1867 107
rect 2000 106 2001 108
rect 2003 106 2004 108
rect 1767 101 1804 102
rect 1526 92 1594 95
rect 1526 90 1528 92
rect 1530 90 1594 92
rect 1526 89 1594 90
rect 1800 91 1804 101
rect 1903 102 1908 103
rect 1903 100 1904 102
rect 1906 100 1908 102
rect 1903 92 1908 100
rect 1800 89 1801 91
rect 1803 89 1804 91
rect 1800 88 1804 89
rect 1817 87 1908 92
rect 928 64 933 79
rect 600 60 933 64
rect 938 73 942 75
rect 938 71 939 73
rect 941 71 942 73
rect 938 63 942 71
rect 938 61 939 63
rect 941 61 942 63
rect 938 60 942 61
rect 952 64 956 79
rect 1080 73 1086 80
rect 1267 79 1348 83
rect 1517 81 1564 85
rect 1817 84 1822 87
rect 1080 71 1082 73
rect 1084 71 1086 73
rect 1080 69 1086 71
rect 1108 73 1113 76
rect 1108 71 1110 73
rect 1112 71 1113 73
rect 952 63 1104 64
rect 952 61 1101 63
rect 1103 61 1104 63
rect 952 60 1104 61
rect 600 56 604 60
rect 1108 56 1113 71
rect 1344 66 1348 79
rect 1344 64 1345 66
rect 1347 64 1348 66
rect 1119 63 1249 64
rect 1119 61 1121 63
rect 1123 62 1249 63
rect 1123 61 1245 62
rect 1119 60 1245 61
rect 1247 60 1249 62
rect 1344 60 1348 64
rect 1358 72 1363 73
rect 1358 70 1360 72
rect 1362 70 1363 72
rect 1240 59 1249 60
rect 1358 56 1363 70
rect 321 55 354 56
rect 321 53 322 55
rect 324 53 349 55
rect 351 53 354 55
rect 321 52 354 53
rect 394 55 459 56
rect 394 53 395 55
rect 397 53 427 55
rect 429 53 454 55
rect 456 53 459 55
rect 394 52 459 53
rect 571 55 604 56
rect 571 53 572 55
rect 574 53 599 55
rect 601 53 604 55
rect 571 52 604 53
rect 644 55 709 56
rect 644 53 645 55
rect 647 53 677 55
rect 679 53 704 55
rect 706 53 709 55
rect 644 52 709 53
rect 821 55 854 56
rect 821 53 822 55
rect 824 53 849 55
rect 851 53 854 55
rect 821 52 854 53
rect 894 55 959 56
rect 894 53 895 55
rect 897 53 927 55
rect 929 53 954 55
rect 956 53 959 55
rect 894 52 959 53
rect 1081 55 1114 56
rect 1081 53 1082 55
rect 1084 53 1109 55
rect 1111 53 1114 55
rect 1081 52 1114 53
rect 1154 55 1219 56
rect 1154 53 1155 55
rect 1157 53 1187 55
rect 1189 53 1214 55
rect 1216 53 1219 55
rect 1154 52 1219 53
rect 1331 55 1364 56
rect 1331 53 1332 55
rect 1334 53 1359 55
rect 1361 53 1364 55
rect 1331 52 1364 53
rect 1404 55 1469 56
rect 1404 53 1405 55
rect 1407 53 1437 55
rect 1439 53 1464 55
rect 1466 53 1469 55
rect 1404 52 1469 53
rect 938 47 942 48
rect 854 45 928 46
rect 854 43 856 45
rect 858 43 928 45
rect 854 42 928 43
rect 61 38 76 39
rect 294 38 325 39
rect 61 36 71 38
rect 73 36 76 38
rect 61 35 76 36
rect 186 37 261 38
rect 186 35 187 37
rect 189 35 258 37
rect 260 35 261 37
rect 294 36 321 38
rect 323 36 325 38
rect 294 35 325 36
rect 438 37 511 38
rect 438 35 439 37
rect 441 35 508 37
rect 510 35 511 37
rect 186 34 261 35
rect 438 34 511 35
rect 688 37 761 38
rect 688 35 689 37
rect 691 35 758 37
rect 760 35 761 37
rect 688 34 761 35
rect 924 31 928 42
rect 938 45 939 47
rect 941 45 942 47
rect 938 38 942 45
rect 938 36 939 38
rect 941 36 942 38
rect 938 35 942 36
rect 954 45 1513 47
rect 954 43 1510 45
rect 1512 43 1513 45
rect 954 42 1513 43
rect 954 31 958 42
rect 1558 39 1564 81
rect 1610 80 1822 84
rect 2000 83 2004 106
rect 1610 56 1614 80
rect 1860 79 2004 83
rect 1800 75 1804 76
rect 1800 73 1801 75
rect 1803 73 1804 75
rect 1581 55 1614 56
rect 1581 53 1582 55
rect 1584 53 1609 55
rect 1611 53 1614 55
rect 1581 52 1614 53
rect 1654 55 1719 56
rect 1654 53 1655 55
rect 1657 53 1687 55
rect 1689 53 1714 55
rect 1716 53 1719 55
rect 1654 52 1719 53
rect 1800 39 1804 73
rect 1860 56 1864 79
rect 1948 73 1952 75
rect 1948 71 1949 73
rect 1951 71 1952 73
rect 1948 63 1952 71
rect 1948 61 1949 63
rect 1951 61 1952 63
rect 1948 60 1952 61
rect 1831 55 1864 56
rect 1831 53 1832 55
rect 1834 53 1859 55
rect 1861 53 1864 55
rect 1831 52 1864 53
rect 1904 55 1969 56
rect 1904 53 1905 55
rect 1907 53 1937 55
rect 1939 53 1964 55
rect 1966 53 1969 55
rect 1904 52 1969 53
rect 1948 47 1952 48
rect 1948 45 1949 47
rect 1951 45 1952 47
rect 1558 38 1591 39
rect 1800 38 1840 39
rect 1080 37 1099 38
rect 1080 35 1082 37
rect 1084 35 1094 37
rect 1096 35 1099 37
rect 1080 34 1099 35
rect 1196 37 1271 38
rect 1196 35 1197 37
rect 1199 35 1268 37
rect 1270 35 1271 37
rect 1196 34 1271 35
rect 1344 37 1348 38
rect 1344 35 1345 37
rect 1347 35 1348 37
rect 1344 34 1348 35
rect 1448 37 1521 38
rect 1448 35 1449 37
rect 1451 35 1518 37
rect 1520 35 1521 37
rect 1558 36 1582 38
rect 1584 36 1591 38
rect 1558 35 1591 36
rect 1698 37 1771 38
rect 1698 35 1699 37
rect 1701 35 1768 37
rect 1770 35 1771 37
rect 1800 36 1832 38
rect 1834 36 1840 38
rect 1800 35 1840 36
rect 1948 38 1952 45
rect 1948 36 1949 38
rect 1951 36 1952 38
rect 1948 35 1952 36
rect 1448 34 1521 35
rect 1698 34 1771 35
rect 39 29 157 30
rect 39 27 40 29
rect 42 27 154 29
rect 156 27 157 29
rect 39 26 157 27
rect 289 29 407 30
rect 289 27 290 29
rect 292 27 404 29
rect 406 27 407 29
rect 289 26 407 27
rect 539 29 657 30
rect 539 27 540 29
rect 542 27 654 29
rect 656 27 657 29
rect 539 26 657 27
rect 789 29 907 30
rect 789 27 790 29
rect 792 27 904 29
rect 906 27 907 29
rect 924 27 958 31
rect 1049 29 1167 30
rect 1049 27 1050 29
rect 1052 27 1164 29
rect 1166 27 1167 29
rect 789 26 907 27
rect 1049 26 1167 27
rect 1299 29 1417 30
rect 1299 27 1300 29
rect 1302 27 1414 29
rect 1416 27 1417 29
rect 1299 26 1417 27
rect 1549 29 1667 30
rect 1549 27 1550 29
rect 1552 27 1664 29
rect 1666 27 1667 29
rect 1549 26 1667 27
rect 1799 29 1917 30
rect 1799 27 1800 29
rect 1802 27 1914 29
rect 1916 27 1917 29
rect 1799 26 1917 27
rect 596 21 600 22
rect 596 19 597 21
rect 599 19 600 21
rect 596 15 600 19
rect 845 21 850 22
rect 845 19 847 21
rect 849 19 850 21
rect 845 4 850 19
rect 29 0 850 4
<< alu3 >>
rect 363 226 1618 233
rect 363 204 368 226
rect 363 202 365 204
rect 367 202 368 204
rect 363 200 368 202
rect 443 221 448 222
rect 443 219 445 221
rect 447 219 448 221
rect 443 200 448 219
rect 568 204 795 209
rect 443 198 444 200
rect 446 198 448 200
rect 443 196 448 198
rect 120 194 124 195
rect 120 192 121 194
rect 123 192 124 194
rect 120 178 124 192
rect 569 186 574 204
rect 569 184 570 186
rect 572 184 574 186
rect 569 178 574 184
rect 120 176 121 178
rect 123 176 124 178
rect 120 175 124 176
rect 124 159 130 160
rect 124 157 126 159
rect 128 157 130 159
rect 113 119 117 121
rect 34 116 38 118
rect 34 114 35 116
rect 37 114 38 116
rect 34 91 38 114
rect 34 89 35 91
rect 37 89 38 91
rect 34 88 38 89
rect 113 117 114 119
rect 116 117 117 119
rect 113 90 117 117
rect 113 88 114 90
rect 116 88 117 90
rect 113 86 117 88
rect 124 4 130 157
rect 655 118 659 119
rect 655 116 656 118
rect 658 116 659 118
rect 655 101 659 116
rect 790 105 795 204
rect 856 208 864 210
rect 856 206 860 208
rect 862 206 864 208
rect 856 128 864 206
rect 873 196 878 200
rect 873 194 875 196
rect 877 194 878 196
rect 873 170 878 194
rect 873 168 874 170
rect 876 168 878 170
rect 873 166 878 168
rect 856 126 858 128
rect 860 126 864 128
rect 856 124 864 126
rect 873 147 878 148
rect 873 145 874 147
rect 876 145 878 147
rect 873 123 878 145
rect 1606 128 1611 226
rect 1606 126 1608 128
rect 1610 126 1611 128
rect 1606 124 1611 126
rect 873 121 874 123
rect 876 121 878 123
rect 873 120 878 121
rect 1017 119 1052 121
rect 1017 117 1018 119
rect 1020 117 1049 119
rect 1051 117 1052 119
rect 1017 116 1052 117
rect 1903 119 1907 120
rect 1903 117 1904 119
rect 1906 117 1907 119
rect 887 105 892 109
rect 790 103 889 105
rect 891 103 892 105
rect 790 101 892 103
rect 1903 102 1907 117
rect 655 99 656 101
rect 658 99 659 101
rect 1903 100 1904 102
rect 1906 100 1907 102
rect 1903 99 1907 100
rect 655 98 659 99
rect 1006 95 1037 97
rect 1006 93 1008 95
rect 1010 93 1032 95
rect 1034 93 1037 95
rect 1006 92 1037 93
rect 1502 92 1533 95
rect 219 91 264 92
rect 219 89 221 91
rect 223 89 256 91
rect 258 89 264 91
rect 219 88 264 89
rect 1255 90 1285 92
rect 1255 88 1257 90
rect 1259 88 1282 90
rect 1284 88 1285 90
rect 1502 90 1503 92
rect 1505 90 1528 92
rect 1530 90 1533 92
rect 1502 89 1533 90
rect 1800 91 1804 92
rect 1800 89 1801 91
rect 1803 89 1804 91
rect 1255 87 1285 88
rect 1080 73 1086 76
rect 1080 71 1082 73
rect 1084 71 1086 73
rect 1800 75 1804 89
rect 1800 73 1801 75
rect 1803 73 1804 75
rect 1800 72 1804 73
rect 938 63 942 64
rect 938 61 939 63
rect 941 61 942 63
rect 938 47 942 61
rect 938 45 939 47
rect 941 45 942 47
rect 938 44 942 45
rect 1080 37 1086 71
rect 1344 66 1348 68
rect 1344 64 1345 66
rect 1347 64 1348 66
rect 1099 63 1125 64
rect 1099 61 1101 63
rect 1103 61 1121 63
rect 1123 61 1125 63
rect 1099 60 1125 61
rect 1080 35 1082 37
rect 1084 35 1086 37
rect 1080 34 1086 35
rect 1344 37 1348 64
rect 1948 63 1952 64
rect 1948 61 1949 63
rect 1951 61 1952 63
rect 1948 47 1952 61
rect 1948 45 1949 47
rect 1951 45 1952 47
rect 1948 44 1952 45
rect 1344 35 1345 37
rect 1347 35 1348 37
rect 1344 33 1348 35
rect 596 21 600 22
rect 596 19 597 21
rect 599 19 600 21
rect 596 4 600 19
rect 124 0 600 4
<< ptie >>
rect 62 226 68 228
rect 62 224 64 226
rect 66 224 68 226
rect 62 222 68 224
rect 102 226 108 228
rect 102 224 104 226
rect 106 224 108 226
rect 102 222 108 224
rect 173 226 179 228
rect 173 224 175 226
rect 177 224 179 226
rect 173 222 179 224
rect 214 226 220 228
rect 214 224 216 226
rect 218 224 220 226
rect 214 222 220 224
rect 364 225 370 227
rect 364 223 366 225
rect 368 223 370 225
rect 364 221 370 223
rect 432 225 438 227
rect 432 223 434 225
rect 436 223 438 225
rect 432 221 438 223
rect 444 225 450 227
rect 444 223 446 225
rect 448 223 450 225
rect 444 221 450 223
rect 485 225 491 227
rect 485 223 487 225
rect 489 223 491 225
rect 485 221 491 223
rect 569 225 575 227
rect 569 223 571 225
rect 573 223 575 225
rect 569 221 575 223
rect 637 225 643 227
rect 637 223 639 225
rect 641 223 643 225
rect 637 221 643 223
rect 649 225 655 227
rect 649 223 651 225
rect 653 223 655 225
rect 649 221 655 223
rect 690 225 696 227
rect 690 223 692 225
rect 694 223 696 225
rect 690 221 696 223
rect 1852 226 1858 228
rect 1852 224 1854 226
rect 1856 224 1858 226
rect 1852 222 1858 224
rect 1892 226 1898 228
rect 1892 224 1894 226
rect 1896 224 1898 226
rect 1892 222 1898 224
rect 1963 226 1969 228
rect 1963 224 1965 226
rect 1967 224 1969 226
rect 1963 222 1969 224
rect 2004 226 2010 228
rect 2004 224 2006 226
rect 2008 224 2010 226
rect 2004 222 2010 224
rect 34 94 40 96
rect 34 92 36 94
rect 38 92 40 94
rect 34 90 40 92
rect 102 94 108 96
rect 102 92 104 94
rect 106 92 108 94
rect 102 90 108 92
rect 114 94 120 96
rect 114 92 116 94
rect 118 92 120 94
rect 114 90 120 92
rect 155 94 161 96
rect 155 92 157 94
rect 159 92 161 94
rect 155 90 161 92
rect 238 94 244 96
rect 238 92 240 94
rect 242 92 244 94
rect 238 90 244 92
rect 279 94 285 96
rect 279 92 281 94
rect 283 92 285 94
rect 279 90 285 92
rect 392 93 398 95
rect 392 91 394 93
rect 396 91 398 93
rect 392 89 398 91
rect 432 93 438 95
rect 432 91 434 93
rect 436 91 438 93
rect 432 89 438 91
rect 503 93 509 95
rect 503 91 505 93
rect 507 91 509 93
rect 503 89 509 91
rect 544 93 550 95
rect 544 91 546 93
rect 548 91 550 93
rect 544 89 550 91
rect 597 93 603 95
rect 597 91 599 93
rect 601 91 603 93
rect 597 89 603 91
rect 637 93 643 95
rect 637 91 639 93
rect 641 91 643 93
rect 637 89 643 91
rect 708 93 714 95
rect 708 91 710 93
rect 712 91 714 93
rect 708 89 714 91
rect 749 93 755 95
rect 749 91 751 93
rect 753 91 755 93
rect 749 89 755 91
rect 776 94 782 96
rect 816 94 822 96
rect 776 92 778 94
rect 780 92 782 94
rect 776 90 782 92
rect 816 92 818 94
rect 820 92 822 94
rect 816 90 822 92
rect 857 94 863 96
rect 857 92 859 94
rect 861 92 863 94
rect 857 90 863 92
rect 921 94 927 96
rect 921 92 923 94
rect 925 92 927 94
rect 921 90 927 92
rect 962 94 968 96
rect 962 92 964 94
rect 966 92 968 94
rect 962 90 968 92
rect 1026 94 1032 96
rect 1066 94 1072 96
rect 1026 92 1028 94
rect 1030 92 1032 94
rect 1026 90 1032 92
rect 1066 92 1068 94
rect 1070 92 1072 94
rect 1066 90 1072 92
rect 1107 94 1113 96
rect 1107 92 1109 94
rect 1111 92 1113 94
rect 1107 90 1113 92
rect 1171 94 1177 96
rect 1171 92 1173 94
rect 1175 92 1177 94
rect 1171 90 1177 92
rect 1212 94 1218 96
rect 1212 92 1214 94
rect 1216 92 1218 94
rect 1212 90 1218 92
rect 1276 94 1282 96
rect 1316 94 1322 96
rect 1276 92 1278 94
rect 1280 92 1282 94
rect 1276 90 1282 92
rect 1316 92 1318 94
rect 1320 92 1322 94
rect 1316 90 1322 92
rect 1357 94 1363 96
rect 1357 92 1359 94
rect 1361 92 1363 94
rect 1357 90 1363 92
rect 1421 94 1427 96
rect 1421 92 1423 94
rect 1425 92 1427 94
rect 1421 90 1427 92
rect 1462 94 1468 96
rect 1462 92 1464 94
rect 1466 92 1468 94
rect 1462 90 1468 92
rect 1526 94 1532 96
rect 1566 94 1572 96
rect 1526 92 1528 94
rect 1530 92 1532 94
rect 1526 90 1532 92
rect 1566 92 1568 94
rect 1570 92 1572 94
rect 1566 90 1572 92
rect 1607 94 1613 96
rect 1607 92 1609 94
rect 1611 92 1613 94
rect 1607 90 1613 92
rect 1671 94 1677 96
rect 1671 92 1673 94
rect 1675 92 1677 94
rect 1671 90 1677 92
rect 1712 94 1718 96
rect 1712 92 1714 94
rect 1716 92 1718 94
rect 1712 90 1718 92
rect 1824 94 1830 96
rect 1824 92 1826 94
rect 1828 92 1830 94
rect 1824 90 1830 92
rect 1892 94 1898 96
rect 1892 92 1894 94
rect 1896 92 1898 94
rect 1892 90 1898 92
rect 1904 94 1910 96
rect 1904 92 1906 94
rect 1908 92 1910 94
rect 1904 90 1910 92
rect 1945 94 1951 96
rect 1945 92 1947 94
rect 1949 92 1951 94
rect 1945 90 1951 92
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 48 72 54 74
rect 48 70 50 72
rect 52 70 54 72
rect 8 68 14 70
rect 48 68 54 70
rect 89 72 95 74
rect 89 70 91 72
rect 93 70 95 72
rect 89 68 95 70
rect 153 72 159 74
rect 153 70 155 72
rect 157 70 159 72
rect 153 68 159 70
rect 194 72 200 74
rect 194 70 196 72
rect 198 70 200 72
rect 194 68 200 70
rect 258 72 264 74
rect 258 70 260 72
rect 262 70 264 72
rect 298 72 304 74
rect 298 70 300 72
rect 302 70 304 72
rect 258 68 264 70
rect 298 68 304 70
rect 339 72 345 74
rect 339 70 341 72
rect 343 70 345 72
rect 339 68 345 70
rect 403 72 409 74
rect 403 70 405 72
rect 407 70 409 72
rect 403 68 409 70
rect 444 72 450 74
rect 444 70 446 72
rect 448 70 450 72
rect 444 68 450 70
rect 508 72 514 74
rect 508 70 510 72
rect 512 70 514 72
rect 548 72 554 74
rect 548 70 550 72
rect 552 70 554 72
rect 508 68 514 70
rect 548 68 554 70
rect 589 72 595 74
rect 589 70 591 72
rect 593 70 595 72
rect 589 68 595 70
rect 653 72 659 74
rect 653 70 655 72
rect 657 70 659 72
rect 653 68 659 70
rect 694 72 700 74
rect 694 70 696 72
rect 698 70 700 72
rect 694 68 700 70
rect 758 72 764 74
rect 758 70 760 72
rect 762 70 764 72
rect 798 72 804 74
rect 798 70 800 72
rect 802 70 804 72
rect 758 68 764 70
rect 798 68 804 70
rect 839 72 845 74
rect 839 70 841 72
rect 843 70 845 72
rect 839 68 845 70
rect 903 72 909 74
rect 903 70 905 72
rect 907 70 909 72
rect 903 68 909 70
rect 944 72 950 74
rect 944 70 946 72
rect 948 70 950 72
rect 944 68 950 70
rect 1018 72 1024 74
rect 1018 70 1020 72
rect 1022 70 1024 72
rect 1058 72 1064 74
rect 1058 70 1060 72
rect 1062 70 1064 72
rect 1018 68 1024 70
rect 1058 68 1064 70
rect 1099 72 1105 74
rect 1099 70 1101 72
rect 1103 70 1105 72
rect 1099 68 1105 70
rect 1163 72 1169 74
rect 1163 70 1165 72
rect 1167 70 1169 72
rect 1163 68 1169 70
rect 1204 72 1210 74
rect 1204 70 1206 72
rect 1208 70 1210 72
rect 1204 68 1210 70
rect 1268 72 1274 74
rect 1268 70 1270 72
rect 1272 70 1274 72
rect 1308 72 1314 74
rect 1308 70 1310 72
rect 1312 70 1314 72
rect 1268 68 1274 70
rect 1308 68 1314 70
rect 1349 72 1355 74
rect 1349 70 1351 72
rect 1353 70 1355 72
rect 1349 68 1355 70
rect 1413 72 1419 74
rect 1413 70 1415 72
rect 1417 70 1419 72
rect 1413 68 1419 70
rect 1454 72 1460 74
rect 1454 70 1456 72
rect 1458 70 1460 72
rect 1454 68 1460 70
rect 1518 72 1524 74
rect 1518 70 1520 72
rect 1522 70 1524 72
rect 1558 72 1564 74
rect 1558 70 1560 72
rect 1562 70 1564 72
rect 1518 68 1524 70
rect 1558 68 1564 70
rect 1599 72 1605 74
rect 1599 70 1601 72
rect 1603 70 1605 72
rect 1599 68 1605 70
rect 1663 72 1669 74
rect 1663 70 1665 72
rect 1667 70 1669 72
rect 1663 68 1669 70
rect 1704 72 1710 74
rect 1704 70 1706 72
rect 1708 70 1710 72
rect 1704 68 1710 70
rect 1768 72 1774 74
rect 1768 70 1770 72
rect 1772 70 1774 72
rect 1808 72 1814 74
rect 1808 70 1810 72
rect 1812 70 1814 72
rect 1768 68 1774 70
rect 1808 68 1814 70
rect 1849 72 1855 74
rect 1849 70 1851 72
rect 1853 70 1855 72
rect 1849 68 1855 70
rect 1913 72 1919 74
rect 1913 70 1915 72
rect 1917 70 1919 72
rect 1913 68 1919 70
rect 1954 72 1960 74
rect 1954 70 1956 72
rect 1958 70 1960 72
rect 1954 68 1960 70
<< ntie >>
rect 62 166 68 168
rect 62 164 64 166
rect 66 164 68 166
rect 62 162 68 164
rect 102 166 108 168
rect 102 164 104 166
rect 106 164 108 166
rect 140 166 146 168
rect 102 162 108 164
rect 140 164 142 166
rect 144 164 146 166
rect 214 166 220 168
rect 140 162 146 164
rect 214 164 216 166
rect 218 164 220 166
rect 214 162 220 164
rect 364 165 370 167
rect 364 163 366 165
rect 368 163 370 165
rect 364 161 370 163
rect 432 165 438 167
rect 432 163 434 165
rect 436 163 438 165
rect 432 161 438 163
rect 444 165 450 167
rect 444 163 446 165
rect 448 163 450 165
rect 518 165 524 167
rect 444 161 450 163
rect 518 163 520 165
rect 522 163 524 165
rect 569 165 575 167
rect 518 161 524 163
rect 569 163 571 165
rect 573 163 575 165
rect 569 161 575 163
rect 637 165 643 167
rect 637 163 639 165
rect 641 163 643 165
rect 637 161 643 163
rect 649 165 655 167
rect 649 163 651 165
rect 653 163 655 165
rect 723 165 729 167
rect 649 161 655 163
rect 723 163 725 165
rect 727 163 729 165
rect 1852 166 1858 168
rect 1852 164 1854 166
rect 1856 164 1858 166
rect 723 161 729 163
rect 1852 162 1858 164
rect 1892 166 1898 168
rect 1892 164 1894 166
rect 1896 164 1898 166
rect 1930 166 1936 168
rect 1892 162 1898 164
rect 1930 164 1932 166
rect 1934 164 1936 166
rect 2004 166 2010 168
rect 1930 162 1936 164
rect 2004 164 2006 166
rect 2008 164 2010 166
rect 2004 162 2010 164
rect 34 154 40 156
rect 34 152 36 154
rect 38 152 40 154
rect 34 150 40 152
rect 102 154 108 156
rect 102 152 104 154
rect 106 152 108 154
rect 102 150 108 152
rect 114 154 120 156
rect 114 152 116 154
rect 118 152 120 154
rect 188 154 194 156
rect 114 150 120 152
rect 188 152 190 154
rect 192 152 194 154
rect 238 154 244 156
rect 188 150 194 152
rect 238 152 240 154
rect 242 152 244 154
rect 312 154 318 156
rect 238 150 244 152
rect 312 152 314 154
rect 316 152 318 154
rect 392 153 398 155
rect 312 150 318 152
rect 392 151 394 153
rect 396 151 398 153
rect 392 149 398 151
rect 432 153 438 155
rect 432 151 434 153
rect 436 151 438 153
rect 470 153 476 155
rect 432 149 438 151
rect 470 151 472 153
rect 474 151 476 153
rect 544 153 550 155
rect 470 149 476 151
rect 544 151 546 153
rect 548 151 550 153
rect 544 149 550 151
rect 597 153 603 155
rect 597 151 599 153
rect 601 151 603 153
rect 597 149 603 151
rect 637 153 643 155
rect 637 151 639 153
rect 641 151 643 153
rect 675 153 681 155
rect 637 149 643 151
rect 675 151 677 153
rect 679 151 681 153
rect 749 153 755 155
rect 675 149 681 151
rect 749 151 751 153
rect 753 151 755 153
rect 749 149 755 151
rect 776 154 782 156
rect 776 152 778 154
rect 780 152 782 154
rect 816 154 822 156
rect 776 150 782 152
rect 816 152 818 154
rect 820 152 822 154
rect 890 154 896 156
rect 816 150 822 152
rect 890 152 892 154
rect 894 152 896 154
rect 921 154 927 156
rect 890 150 896 152
rect 921 152 923 154
rect 925 152 927 154
rect 995 154 1001 156
rect 921 150 927 152
rect 995 152 997 154
rect 999 152 1001 154
rect 1026 154 1032 156
rect 995 150 1001 152
rect 1026 152 1028 154
rect 1030 152 1032 154
rect 1066 154 1072 156
rect 1026 150 1032 152
rect 1066 152 1068 154
rect 1070 152 1072 154
rect 1140 154 1146 156
rect 1066 150 1072 152
rect 1140 152 1142 154
rect 1144 152 1146 154
rect 1171 154 1177 156
rect 1140 150 1146 152
rect 1171 152 1173 154
rect 1175 152 1177 154
rect 1245 154 1251 156
rect 1171 150 1177 152
rect 1245 152 1247 154
rect 1249 152 1251 154
rect 1276 154 1282 156
rect 1245 150 1251 152
rect 1276 152 1278 154
rect 1280 152 1282 154
rect 1316 154 1322 156
rect 1276 150 1282 152
rect 1316 152 1318 154
rect 1320 152 1322 154
rect 1390 154 1396 156
rect 1316 150 1322 152
rect 1390 152 1392 154
rect 1394 152 1396 154
rect 1421 154 1427 156
rect 1390 150 1396 152
rect 1421 152 1423 154
rect 1425 152 1427 154
rect 1495 154 1501 156
rect 1421 150 1427 152
rect 1495 152 1497 154
rect 1499 152 1501 154
rect 1526 154 1532 156
rect 1495 150 1501 152
rect 1526 152 1528 154
rect 1530 152 1532 154
rect 1566 154 1572 156
rect 1526 150 1532 152
rect 1566 152 1568 154
rect 1570 152 1572 154
rect 1640 154 1646 156
rect 1566 150 1572 152
rect 1640 152 1642 154
rect 1644 152 1646 154
rect 1671 154 1677 156
rect 1640 150 1646 152
rect 1671 152 1673 154
rect 1675 152 1677 154
rect 1745 154 1751 156
rect 1671 150 1677 152
rect 1745 152 1747 154
rect 1749 152 1751 154
rect 1824 154 1830 156
rect 1745 150 1751 152
rect 1824 152 1826 154
rect 1828 152 1830 154
rect 1824 150 1830 152
rect 1892 154 1898 156
rect 1892 152 1894 154
rect 1896 152 1898 154
rect 1892 150 1898 152
rect 1904 154 1910 156
rect 1904 152 1906 154
rect 1908 152 1910 154
rect 1978 154 1984 156
rect 1904 150 1910 152
rect 1978 152 1980 154
rect 1982 152 1984 154
rect 1978 150 1984 152
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 48 12 54 14
rect 8 8 14 10
rect 48 10 50 12
rect 52 10 54 12
rect 122 12 128 14
rect 48 8 54 10
rect 122 10 124 12
rect 126 10 128 12
rect 153 12 159 14
rect 122 8 128 10
rect 153 10 155 12
rect 157 10 159 12
rect 227 12 233 14
rect 153 8 159 10
rect 227 10 229 12
rect 231 10 233 12
rect 258 12 264 14
rect 227 8 233 10
rect 258 10 260 12
rect 262 10 264 12
rect 298 12 304 14
rect 258 8 264 10
rect 298 10 300 12
rect 302 10 304 12
rect 372 12 378 14
rect 298 8 304 10
rect 372 10 374 12
rect 376 10 378 12
rect 403 12 409 14
rect 372 8 378 10
rect 403 10 405 12
rect 407 10 409 12
rect 477 12 483 14
rect 403 8 409 10
rect 477 10 479 12
rect 481 10 483 12
rect 508 12 514 14
rect 477 8 483 10
rect 508 10 510 12
rect 512 10 514 12
rect 548 12 554 14
rect 508 8 514 10
rect 548 10 550 12
rect 552 10 554 12
rect 622 12 628 14
rect 548 8 554 10
rect 622 10 624 12
rect 626 10 628 12
rect 653 12 659 14
rect 622 8 628 10
rect 653 10 655 12
rect 657 10 659 12
rect 727 12 733 14
rect 653 8 659 10
rect 727 10 729 12
rect 731 10 733 12
rect 758 12 764 14
rect 727 8 733 10
rect 758 10 760 12
rect 762 10 764 12
rect 798 12 804 14
rect 758 8 764 10
rect 798 10 800 12
rect 802 10 804 12
rect 872 12 878 14
rect 798 8 804 10
rect 872 10 874 12
rect 876 10 878 12
rect 903 12 909 14
rect 872 8 878 10
rect 903 10 905 12
rect 907 10 909 12
rect 977 12 983 14
rect 903 8 909 10
rect 977 10 979 12
rect 981 10 983 12
rect 1018 12 1024 14
rect 977 8 983 10
rect 1018 10 1020 12
rect 1022 10 1024 12
rect 1058 12 1064 14
rect 1018 8 1024 10
rect 1058 10 1060 12
rect 1062 10 1064 12
rect 1132 12 1138 14
rect 1058 8 1064 10
rect 1132 10 1134 12
rect 1136 10 1138 12
rect 1163 12 1169 14
rect 1132 8 1138 10
rect 1163 10 1165 12
rect 1167 10 1169 12
rect 1237 12 1243 14
rect 1163 8 1169 10
rect 1237 10 1239 12
rect 1241 10 1243 12
rect 1268 12 1274 14
rect 1237 8 1243 10
rect 1268 10 1270 12
rect 1272 10 1274 12
rect 1308 12 1314 14
rect 1268 8 1274 10
rect 1308 10 1310 12
rect 1312 10 1314 12
rect 1382 12 1388 14
rect 1308 8 1314 10
rect 1382 10 1384 12
rect 1386 10 1388 12
rect 1413 12 1419 14
rect 1382 8 1388 10
rect 1413 10 1415 12
rect 1417 10 1419 12
rect 1487 12 1493 14
rect 1413 8 1419 10
rect 1487 10 1489 12
rect 1491 10 1493 12
rect 1518 12 1524 14
rect 1487 8 1493 10
rect 1518 10 1520 12
rect 1522 10 1524 12
rect 1558 12 1564 14
rect 1518 8 1524 10
rect 1558 10 1560 12
rect 1562 10 1564 12
rect 1632 12 1638 14
rect 1558 8 1564 10
rect 1632 10 1634 12
rect 1636 10 1638 12
rect 1663 12 1669 14
rect 1632 8 1638 10
rect 1663 10 1665 12
rect 1667 10 1669 12
rect 1737 12 1743 14
rect 1663 8 1669 10
rect 1737 10 1739 12
rect 1741 10 1743 12
rect 1768 12 1774 14
rect 1737 8 1743 10
rect 1768 10 1770 12
rect 1772 10 1774 12
rect 1808 12 1814 14
rect 1768 8 1774 10
rect 1808 10 1810 12
rect 1812 10 1814 12
rect 1882 12 1888 14
rect 1808 8 1814 10
rect 1882 10 1884 12
rect 1886 10 1888 12
rect 1913 12 1919 14
rect 1882 8 1888 10
rect 1913 10 1915 12
rect 1917 10 1919 12
rect 1987 12 1993 14
rect 1913 8 1919 10
rect 1987 10 1989 12
rect 1991 10 1993 12
rect 1987 8 1993 10
<< nmos >>
rect 40 207 42 218
rect 47 207 49 218
rect 60 207 62 216
rect 80 207 82 218
rect 87 207 89 218
rect 100 207 102 216
rect 128 210 130 222
rect 135 210 137 222
rect 145 210 147 219
rect 155 210 157 219
rect 171 205 173 214
rect 192 207 194 218
rect 199 207 201 218
rect 212 207 214 216
rect 370 206 372 215
rect 383 206 385 217
rect 390 206 392 217
rect 410 206 412 217
rect 417 206 419 217
rect 430 206 432 215
rect 450 206 452 215
rect 463 206 465 217
rect 470 206 472 217
rect 491 204 493 213
rect 507 209 509 218
rect 517 209 519 218
rect 527 209 529 221
rect 534 209 536 221
rect 575 206 577 215
rect 588 206 590 217
rect 595 206 597 217
rect 615 206 617 217
rect 622 206 624 217
rect 635 206 637 215
rect 655 206 657 215
rect 668 206 670 217
rect 675 206 677 217
rect 696 204 698 213
rect 712 209 714 218
rect 722 209 724 218
rect 732 209 734 221
rect 739 209 741 221
rect 1830 207 1832 218
rect 1837 207 1839 218
rect 1850 207 1852 216
rect 1870 207 1872 218
rect 1877 207 1879 218
rect 1890 207 1892 216
rect 1918 210 1920 222
rect 1925 210 1927 222
rect 1935 210 1937 219
rect 1945 210 1947 219
rect 1961 205 1963 214
rect 1982 207 1984 218
rect 1989 207 1991 218
rect 2002 207 2004 216
rect 40 102 42 111
rect 53 100 55 111
rect 60 100 62 111
rect 80 100 82 111
rect 87 100 89 111
rect 100 102 102 111
rect 120 102 122 111
rect 133 100 135 111
rect 140 100 142 111
rect 161 104 163 113
rect 177 99 179 108
rect 187 99 189 108
rect 197 96 199 108
rect 204 96 206 108
rect 244 102 246 111
rect 257 100 259 111
rect 264 100 266 111
rect 285 104 287 113
rect 301 99 303 108
rect 311 99 313 108
rect 321 96 323 108
rect 328 96 330 108
rect 370 99 372 110
rect 377 99 379 110
rect 390 101 392 110
rect 410 99 412 110
rect 417 99 419 110
rect 430 101 432 110
rect 458 95 460 107
rect 465 95 467 107
rect 475 98 477 107
rect 485 98 487 107
rect 501 103 503 112
rect 522 99 524 110
rect 529 99 531 110
rect 542 101 544 110
rect 575 99 577 110
rect 582 99 584 110
rect 595 101 597 110
rect 615 99 617 110
rect 622 99 624 110
rect 635 101 637 110
rect 663 95 665 107
rect 670 95 672 107
rect 680 98 682 107
rect 690 98 692 107
rect 706 103 708 112
rect 727 99 729 110
rect 734 99 736 110
rect 747 101 749 110
rect 782 104 784 113
rect 792 107 794 113
rect 802 107 804 113
rect 822 102 824 111
rect 835 100 837 111
rect 842 100 844 111
rect 863 104 865 113
rect 879 99 881 108
rect 889 99 891 108
rect 899 96 901 108
rect 906 96 908 108
rect 927 102 929 111
rect 940 100 942 111
rect 947 100 949 111
rect 968 104 970 113
rect 984 99 986 108
rect 994 99 996 108
rect 1004 96 1006 108
rect 1011 96 1013 108
rect 1032 104 1034 113
rect 1042 107 1044 113
rect 1052 107 1054 113
rect 1072 102 1074 111
rect 1085 100 1087 111
rect 1092 100 1094 111
rect 1113 104 1115 113
rect 1129 99 1131 108
rect 1139 99 1141 108
rect 1149 96 1151 108
rect 1156 96 1158 108
rect 1177 102 1179 111
rect 1190 100 1192 111
rect 1197 100 1199 111
rect 1218 104 1220 113
rect 1234 99 1236 108
rect 1244 99 1246 108
rect 1254 96 1256 108
rect 1261 96 1263 108
rect 1282 104 1284 113
rect 1292 107 1294 113
rect 1302 107 1304 113
rect 1322 102 1324 111
rect 1335 100 1337 111
rect 1342 100 1344 111
rect 1363 104 1365 113
rect 1379 99 1381 108
rect 1389 99 1391 108
rect 1399 96 1401 108
rect 1406 96 1408 108
rect 1427 102 1429 111
rect 1440 100 1442 111
rect 1447 100 1449 111
rect 1468 104 1470 113
rect 1484 99 1486 108
rect 1494 99 1496 108
rect 1504 96 1506 108
rect 1511 96 1513 108
rect 1532 104 1534 113
rect 1542 107 1544 113
rect 1552 107 1554 113
rect 1572 102 1574 111
rect 1585 100 1587 111
rect 1592 100 1594 111
rect 1613 104 1615 113
rect 1629 99 1631 108
rect 1639 99 1641 108
rect 1649 96 1651 108
rect 1656 96 1658 108
rect 1677 102 1679 111
rect 1690 100 1692 111
rect 1697 100 1699 111
rect 1718 104 1720 113
rect 1734 99 1736 108
rect 1744 99 1746 108
rect 1754 96 1756 108
rect 1761 96 1763 108
rect 1830 102 1832 111
rect 1843 100 1845 111
rect 1850 100 1852 111
rect 1870 100 1872 111
rect 1877 100 1879 111
rect 1890 102 1892 111
rect 1910 102 1912 111
rect 1923 100 1925 111
rect 1930 100 1932 111
rect 1951 104 1953 113
rect 1967 99 1969 108
rect 1977 99 1979 108
rect 1987 96 1989 108
rect 1994 96 1996 108
rect 14 51 16 60
rect 24 51 26 57
rect 34 51 36 57
rect 54 53 56 62
rect 67 53 69 64
rect 74 53 76 64
rect 95 51 97 60
rect 111 56 113 65
rect 121 56 123 65
rect 131 56 133 68
rect 138 56 140 68
rect 159 53 161 62
rect 172 53 174 64
rect 179 53 181 64
rect 200 51 202 60
rect 216 56 218 65
rect 226 56 228 65
rect 236 56 238 68
rect 243 56 245 68
rect 264 51 266 60
rect 274 51 276 57
rect 284 51 286 57
rect 304 53 306 62
rect 317 53 319 64
rect 324 53 326 64
rect 345 51 347 60
rect 361 56 363 65
rect 371 56 373 65
rect 381 56 383 68
rect 388 56 390 68
rect 409 53 411 62
rect 422 53 424 64
rect 429 53 431 64
rect 450 51 452 60
rect 466 56 468 65
rect 476 56 478 65
rect 486 56 488 68
rect 493 56 495 68
rect 514 51 516 60
rect 524 51 526 57
rect 534 51 536 57
rect 554 53 556 62
rect 567 53 569 64
rect 574 53 576 64
rect 595 51 597 60
rect 611 56 613 65
rect 621 56 623 65
rect 631 56 633 68
rect 638 56 640 68
rect 659 53 661 62
rect 672 53 674 64
rect 679 53 681 64
rect 700 51 702 60
rect 716 56 718 65
rect 726 56 728 65
rect 736 56 738 68
rect 743 56 745 68
rect 764 51 766 60
rect 774 51 776 57
rect 784 51 786 57
rect 804 53 806 62
rect 817 53 819 64
rect 824 53 826 64
rect 845 51 847 60
rect 861 56 863 65
rect 871 56 873 65
rect 881 56 883 68
rect 888 56 890 68
rect 909 53 911 62
rect 922 53 924 64
rect 929 53 931 64
rect 950 51 952 60
rect 966 56 968 65
rect 976 56 978 65
rect 986 56 988 68
rect 993 56 995 68
rect 1024 51 1026 60
rect 1034 51 1036 57
rect 1044 51 1046 57
rect 1064 53 1066 62
rect 1077 53 1079 64
rect 1084 53 1086 64
rect 1105 51 1107 60
rect 1121 56 1123 65
rect 1131 56 1133 65
rect 1141 56 1143 68
rect 1148 56 1150 68
rect 1169 53 1171 62
rect 1182 53 1184 64
rect 1189 53 1191 64
rect 1210 51 1212 60
rect 1226 56 1228 65
rect 1236 56 1238 65
rect 1246 56 1248 68
rect 1253 56 1255 68
rect 1274 51 1276 60
rect 1284 51 1286 57
rect 1294 51 1296 57
rect 1314 53 1316 62
rect 1327 53 1329 64
rect 1334 53 1336 64
rect 1355 51 1357 60
rect 1371 56 1373 65
rect 1381 56 1383 65
rect 1391 56 1393 68
rect 1398 56 1400 68
rect 1419 53 1421 62
rect 1432 53 1434 64
rect 1439 53 1441 64
rect 1460 51 1462 60
rect 1476 56 1478 65
rect 1486 56 1488 65
rect 1496 56 1498 68
rect 1503 56 1505 68
rect 1524 51 1526 60
rect 1534 51 1536 57
rect 1544 51 1546 57
rect 1564 53 1566 62
rect 1577 53 1579 64
rect 1584 53 1586 64
rect 1605 51 1607 60
rect 1621 56 1623 65
rect 1631 56 1633 65
rect 1641 56 1643 68
rect 1648 56 1650 68
rect 1669 53 1671 62
rect 1682 53 1684 64
rect 1689 53 1691 64
rect 1710 51 1712 60
rect 1726 56 1728 65
rect 1736 56 1738 65
rect 1746 56 1748 68
rect 1753 56 1755 68
rect 1774 51 1776 60
rect 1784 51 1786 57
rect 1794 51 1796 57
rect 1814 53 1816 62
rect 1827 53 1829 64
rect 1834 53 1836 64
rect 1855 51 1857 60
rect 1871 56 1873 65
rect 1881 56 1883 65
rect 1891 56 1893 68
rect 1898 56 1900 68
rect 1919 53 1921 62
rect 1932 53 1934 64
rect 1939 53 1941 64
rect 1960 51 1962 60
rect 1976 56 1978 65
rect 1986 56 1988 65
rect 1996 56 1998 68
rect 2003 56 2005 68
<< pmos >>
rect 40 172 42 185
rect 50 172 52 185
rect 60 174 62 192
rect 80 172 82 185
rect 90 172 92 185
rect 100 174 102 192
rect 127 165 129 192
rect 137 174 139 192
rect 147 174 149 192
rect 163 165 165 192
rect 192 172 194 185
rect 202 172 204 185
rect 212 174 214 192
rect 370 173 372 191
rect 380 171 382 184
rect 390 171 392 184
rect 410 171 412 184
rect 420 171 422 184
rect 430 173 432 191
rect 450 173 452 191
rect 460 171 462 184
rect 470 171 472 184
rect 499 164 501 191
rect 515 173 517 191
rect 525 173 527 191
rect 535 164 537 191
rect 575 173 577 191
rect 585 171 587 184
rect 595 171 597 184
rect 615 171 617 184
rect 625 171 627 184
rect 635 173 637 191
rect 655 173 657 191
rect 665 171 667 184
rect 675 171 677 184
rect 704 164 706 191
rect 720 173 722 191
rect 730 173 732 191
rect 740 164 742 191
rect 1830 172 1832 185
rect 1840 172 1842 185
rect 1850 174 1852 192
rect 1870 172 1872 185
rect 1880 172 1882 185
rect 1890 174 1892 192
rect 1917 165 1919 192
rect 1927 174 1929 192
rect 1937 174 1939 192
rect 1953 165 1955 192
rect 1982 172 1984 185
rect 1992 172 1994 185
rect 2002 174 2004 192
rect 40 126 42 144
rect 50 133 52 146
rect 60 133 62 146
rect 80 133 82 146
rect 90 133 92 146
rect 100 126 102 144
rect 120 126 122 144
rect 130 133 132 146
rect 140 133 142 146
rect 169 126 171 153
rect 185 126 187 144
rect 195 126 197 144
rect 205 126 207 153
rect 244 126 246 144
rect 254 133 256 146
rect 264 133 266 146
rect 293 126 295 153
rect 309 126 311 144
rect 319 126 321 144
rect 329 126 331 153
rect 370 132 372 145
rect 380 132 382 145
rect 390 125 392 143
rect 410 132 412 145
rect 420 132 422 145
rect 430 125 432 143
rect 457 125 459 152
rect 467 125 469 143
rect 477 125 479 143
rect 493 125 495 152
rect 522 132 524 145
rect 532 132 534 145
rect 542 125 544 143
rect 575 132 577 145
rect 585 132 587 145
rect 595 125 597 143
rect 615 132 617 145
rect 625 132 627 145
rect 635 125 637 143
rect 662 125 664 152
rect 672 125 674 143
rect 682 125 684 143
rect 698 125 700 152
rect 727 132 729 145
rect 737 132 739 145
rect 747 125 749 143
rect 782 125 784 143
rect 795 132 797 153
rect 802 132 804 153
rect 822 126 824 144
rect 832 133 834 146
rect 842 133 844 146
rect 871 126 873 153
rect 887 126 889 144
rect 897 126 899 144
rect 907 126 909 153
rect 927 126 929 144
rect 937 133 939 146
rect 947 133 949 146
rect 976 126 978 153
rect 992 126 994 144
rect 1002 126 1004 144
rect 1012 126 1014 153
rect 1032 125 1034 143
rect 1045 132 1047 153
rect 1052 132 1054 153
rect 1072 126 1074 144
rect 1082 133 1084 146
rect 1092 133 1094 146
rect 1121 126 1123 153
rect 1137 126 1139 144
rect 1147 126 1149 144
rect 1157 126 1159 153
rect 1177 126 1179 144
rect 1187 133 1189 146
rect 1197 133 1199 146
rect 1226 126 1228 153
rect 1242 126 1244 144
rect 1252 126 1254 144
rect 1262 126 1264 153
rect 1282 125 1284 143
rect 1295 132 1297 153
rect 1302 132 1304 153
rect 1322 126 1324 144
rect 1332 133 1334 146
rect 1342 133 1344 146
rect 1371 126 1373 153
rect 1387 126 1389 144
rect 1397 126 1399 144
rect 1407 126 1409 153
rect 1427 126 1429 144
rect 1437 133 1439 146
rect 1447 133 1449 146
rect 1476 126 1478 153
rect 1492 126 1494 144
rect 1502 126 1504 144
rect 1512 126 1514 153
rect 1532 125 1534 143
rect 1545 132 1547 153
rect 1552 132 1554 153
rect 1572 126 1574 144
rect 1582 133 1584 146
rect 1592 133 1594 146
rect 1621 126 1623 153
rect 1637 126 1639 144
rect 1647 126 1649 144
rect 1657 126 1659 153
rect 1677 126 1679 144
rect 1687 133 1689 146
rect 1697 133 1699 146
rect 1726 126 1728 153
rect 1742 126 1744 144
rect 1752 126 1754 144
rect 1762 126 1764 153
rect 1830 126 1832 144
rect 1840 133 1842 146
rect 1850 133 1852 146
rect 1870 133 1872 146
rect 1880 133 1882 146
rect 1890 126 1892 144
rect 1910 126 1912 144
rect 1920 133 1922 146
rect 1930 133 1932 146
rect 1959 126 1961 153
rect 1975 126 1977 144
rect 1985 126 1987 144
rect 1995 126 1997 153
rect 14 21 16 39
rect 27 11 29 32
rect 34 11 36 32
rect 54 20 56 38
rect 64 18 66 31
rect 74 18 76 31
rect 103 11 105 38
rect 119 20 121 38
rect 129 20 131 38
rect 139 11 141 38
rect 159 20 161 38
rect 169 18 171 31
rect 179 18 181 31
rect 208 11 210 38
rect 224 20 226 38
rect 234 20 236 38
rect 244 11 246 38
rect 264 21 266 39
rect 277 11 279 32
rect 284 11 286 32
rect 304 20 306 38
rect 314 18 316 31
rect 324 18 326 31
rect 353 11 355 38
rect 369 20 371 38
rect 379 20 381 38
rect 389 11 391 38
rect 409 20 411 38
rect 419 18 421 31
rect 429 18 431 31
rect 458 11 460 38
rect 474 20 476 38
rect 484 20 486 38
rect 494 11 496 38
rect 514 21 516 39
rect 527 11 529 32
rect 534 11 536 32
rect 554 20 556 38
rect 564 18 566 31
rect 574 18 576 31
rect 603 11 605 38
rect 619 20 621 38
rect 629 20 631 38
rect 639 11 641 38
rect 659 20 661 38
rect 669 18 671 31
rect 679 18 681 31
rect 708 11 710 38
rect 724 20 726 38
rect 734 20 736 38
rect 744 11 746 38
rect 764 21 766 39
rect 777 11 779 32
rect 784 11 786 32
rect 804 20 806 38
rect 814 18 816 31
rect 824 18 826 31
rect 853 11 855 38
rect 869 20 871 38
rect 879 20 881 38
rect 889 11 891 38
rect 909 20 911 38
rect 919 18 921 31
rect 929 18 931 31
rect 958 11 960 38
rect 974 20 976 38
rect 984 20 986 38
rect 994 11 996 38
rect 1024 21 1026 39
rect 1037 11 1039 32
rect 1044 11 1046 32
rect 1064 20 1066 38
rect 1074 18 1076 31
rect 1084 18 1086 31
rect 1113 11 1115 38
rect 1129 20 1131 38
rect 1139 20 1141 38
rect 1149 11 1151 38
rect 1169 20 1171 38
rect 1179 18 1181 31
rect 1189 18 1191 31
rect 1218 11 1220 38
rect 1234 20 1236 38
rect 1244 20 1246 38
rect 1254 11 1256 38
rect 1274 21 1276 39
rect 1287 11 1289 32
rect 1294 11 1296 32
rect 1314 20 1316 38
rect 1324 18 1326 31
rect 1334 18 1336 31
rect 1363 11 1365 38
rect 1379 20 1381 38
rect 1389 20 1391 38
rect 1399 11 1401 38
rect 1419 20 1421 38
rect 1429 18 1431 31
rect 1439 18 1441 31
rect 1468 11 1470 38
rect 1484 20 1486 38
rect 1494 20 1496 38
rect 1504 11 1506 38
rect 1524 21 1526 39
rect 1537 11 1539 32
rect 1544 11 1546 32
rect 1564 20 1566 38
rect 1574 18 1576 31
rect 1584 18 1586 31
rect 1613 11 1615 38
rect 1629 20 1631 38
rect 1639 20 1641 38
rect 1649 11 1651 38
rect 1669 20 1671 38
rect 1679 18 1681 31
rect 1689 18 1691 31
rect 1718 11 1720 38
rect 1734 20 1736 38
rect 1744 20 1746 38
rect 1754 11 1756 38
rect 1774 21 1776 39
rect 1787 11 1789 32
rect 1794 11 1796 32
rect 1814 20 1816 38
rect 1824 18 1826 31
rect 1834 18 1836 31
rect 1863 11 1865 38
rect 1879 20 1881 38
rect 1889 20 1891 38
rect 1899 11 1901 38
rect 1919 20 1921 38
rect 1929 18 1931 31
rect 1939 18 1941 31
rect 1968 11 1970 38
rect 1984 20 1986 38
rect 1994 20 1996 38
rect 2004 11 2006 38
<< polyct0 >>
rect 58 198 60 200
rect 98 198 100 200
rect 129 197 131 199
rect 139 198 141 200
rect 210 198 212 200
rect 372 197 374 199
rect 428 197 430 199
rect 452 197 454 199
rect 523 197 525 199
rect 533 196 535 198
rect 577 197 579 199
rect 633 197 635 199
rect 657 197 659 199
rect 728 197 730 199
rect 738 196 740 198
rect 1848 198 1850 200
rect 1888 198 1890 200
rect 1919 197 1921 199
rect 1929 198 1931 200
rect 2000 198 2002 200
rect 42 118 44 120
rect 98 118 100 120
rect 122 118 124 120
rect 193 118 195 120
rect 203 119 205 121
rect 246 118 248 120
rect 317 118 319 120
rect 327 119 329 121
rect 388 117 390 119
rect 428 117 430 119
rect 459 118 461 120
rect 469 117 471 119
rect 540 117 542 119
rect 593 117 595 119
rect 633 117 635 119
rect 664 118 666 120
rect 674 117 676 119
rect 745 117 747 119
rect 784 118 786 120
rect 824 118 826 120
rect 895 118 897 120
rect 905 119 907 121
rect 929 118 931 120
rect 1000 118 1002 120
rect 1010 119 1012 121
rect 1034 118 1036 120
rect 1074 118 1076 120
rect 1145 118 1147 120
rect 1155 119 1157 121
rect 1179 118 1181 120
rect 1250 118 1252 120
rect 1260 119 1262 121
rect 1284 118 1286 120
rect 1324 118 1326 120
rect 1395 118 1397 120
rect 1405 119 1407 121
rect 1429 118 1431 120
rect 1500 118 1502 120
rect 1510 119 1512 121
rect 1534 118 1536 120
rect 1574 118 1576 120
rect 1645 118 1647 120
rect 1655 119 1657 121
rect 1679 118 1681 120
rect 1750 118 1752 120
rect 1760 119 1762 121
rect 1832 118 1834 120
rect 1888 118 1890 120
rect 1912 118 1914 120
rect 1983 118 1985 120
rect 1993 119 1995 121
rect 16 44 18 46
rect 56 44 58 46
rect 127 44 129 46
rect 137 43 139 45
rect 161 44 163 46
rect 232 44 234 46
rect 242 43 244 45
rect 266 44 268 46
rect 306 44 308 46
rect 377 44 379 46
rect 387 43 389 45
rect 411 44 413 46
rect 482 44 484 46
rect 492 43 494 45
rect 516 44 518 46
rect 556 44 558 46
rect 627 44 629 46
rect 637 43 639 45
rect 661 44 663 46
rect 732 44 734 46
rect 742 43 744 45
rect 766 44 768 46
rect 806 44 808 46
rect 877 44 879 46
rect 887 43 889 45
rect 911 44 913 46
rect 982 44 984 46
rect 992 43 994 45
rect 1026 44 1028 46
rect 1066 44 1068 46
rect 1137 44 1139 46
rect 1147 43 1149 45
rect 1171 44 1173 46
rect 1242 44 1244 46
rect 1252 43 1254 45
rect 1276 44 1278 46
rect 1316 44 1318 46
rect 1387 44 1389 46
rect 1397 43 1399 45
rect 1421 44 1423 46
rect 1492 44 1494 46
rect 1502 43 1504 45
rect 1526 44 1528 46
rect 1566 44 1568 46
rect 1637 44 1639 46
rect 1647 43 1649 45
rect 1671 44 1673 46
rect 1742 44 1744 46
rect 1752 43 1754 45
rect 1776 44 1778 46
rect 1816 44 1818 46
rect 1887 44 1889 46
rect 1897 43 1899 45
rect 1921 44 1923 46
rect 1992 44 1994 46
rect 2002 43 2004 45
<< polyct1 >>
rect 48 198 50 200
rect 38 190 40 192
rect 88 198 90 200
rect 160 203 162 205
rect 78 190 80 192
rect 200 198 202 200
rect 176 190 178 192
rect 190 190 192 192
rect 382 197 384 199
rect 418 197 420 199
rect 392 189 394 191
rect 408 189 410 191
rect 462 197 464 199
rect 502 202 504 204
rect 472 189 474 191
rect 587 197 589 199
rect 486 189 488 191
rect 623 197 625 199
rect 597 189 599 191
rect 613 189 615 191
rect 667 197 669 199
rect 707 202 709 204
rect 677 189 679 191
rect 1838 198 1840 200
rect 691 189 693 191
rect 1828 190 1830 192
rect 1878 198 1880 200
rect 1950 203 1952 205
rect 1868 190 1870 192
rect 1990 198 1992 200
rect 1966 190 1968 192
rect 1980 190 1982 192
rect 62 126 64 128
rect 78 126 80 128
rect 52 118 54 120
rect 88 118 90 120
rect 142 126 144 128
rect 156 126 158 128
rect 132 118 134 120
rect 266 126 268 128
rect 280 126 282 128
rect 172 113 174 115
rect 256 118 258 120
rect 368 125 370 127
rect 296 113 298 115
rect 408 125 410 127
rect 378 117 380 119
rect 506 125 508 127
rect 418 117 420 119
rect 520 125 522 127
rect 490 112 492 114
rect 573 125 575 127
rect 530 117 532 119
rect 613 125 615 127
rect 583 117 585 119
rect 711 125 713 127
rect 623 117 625 119
rect 725 125 727 127
rect 695 112 697 114
rect 735 117 737 119
rect 804 125 806 127
rect 794 118 796 120
rect 844 126 846 128
rect 858 126 860 128
rect 834 118 836 120
rect 949 126 951 128
rect 963 126 965 128
rect 874 113 876 115
rect 939 118 941 120
rect 1054 125 1056 127
rect 979 113 981 115
rect 1044 118 1046 120
rect 1094 126 1096 128
rect 1108 126 1110 128
rect 1084 118 1086 120
rect 1199 126 1201 128
rect 1213 126 1215 128
rect 1124 113 1126 115
rect 1189 118 1191 120
rect 1304 125 1306 127
rect 1229 113 1231 115
rect 1294 118 1296 120
rect 1344 126 1346 128
rect 1358 126 1360 128
rect 1334 118 1336 120
rect 1449 126 1451 128
rect 1463 126 1465 128
rect 1374 113 1376 115
rect 1439 118 1441 120
rect 1554 125 1556 127
rect 1479 113 1481 115
rect 1544 118 1546 120
rect 1594 126 1596 128
rect 1608 126 1610 128
rect 1584 118 1586 120
rect 1699 126 1701 128
rect 1713 126 1715 128
rect 1624 113 1626 115
rect 1689 118 1691 120
rect 1852 126 1854 128
rect 1868 126 1870 128
rect 1729 113 1731 115
rect 1842 118 1844 120
rect 1878 118 1880 120
rect 1932 126 1934 128
rect 1946 126 1948 128
rect 1922 118 1924 120
rect 1962 113 1964 115
rect 26 44 28 46
rect 66 44 68 46
rect 36 37 38 39
rect 106 49 108 51
rect 76 36 78 38
rect 171 44 173 46
rect 90 36 92 38
rect 211 49 213 51
rect 181 36 183 38
rect 276 44 278 46
rect 195 36 197 38
rect 316 44 318 46
rect 286 37 288 39
rect 356 49 358 51
rect 326 36 328 38
rect 421 44 423 46
rect 340 36 342 38
rect 461 49 463 51
rect 431 36 433 38
rect 526 44 528 46
rect 445 36 447 38
rect 566 44 568 46
rect 536 37 538 39
rect 606 49 608 51
rect 576 36 578 38
rect 671 44 673 46
rect 590 36 592 38
rect 711 49 713 51
rect 681 36 683 38
rect 776 44 778 46
rect 695 36 697 38
rect 816 44 818 46
rect 786 37 788 39
rect 856 49 858 51
rect 826 36 828 38
rect 921 44 923 46
rect 840 36 842 38
rect 961 49 963 51
rect 931 36 933 38
rect 1036 44 1038 46
rect 945 36 947 38
rect 1076 44 1078 46
rect 1046 37 1048 39
rect 1116 49 1118 51
rect 1086 36 1088 38
rect 1181 44 1183 46
rect 1100 36 1102 38
rect 1221 49 1223 51
rect 1191 36 1193 38
rect 1286 44 1288 46
rect 1205 36 1207 38
rect 1326 44 1328 46
rect 1296 37 1298 39
rect 1366 49 1368 51
rect 1336 36 1338 38
rect 1431 44 1433 46
rect 1350 36 1352 38
rect 1471 49 1473 51
rect 1441 36 1443 38
rect 1536 44 1538 46
rect 1455 36 1457 38
rect 1576 44 1578 46
rect 1546 37 1548 39
rect 1616 49 1618 51
rect 1586 36 1588 38
rect 1681 44 1683 46
rect 1600 36 1602 38
rect 1721 49 1723 51
rect 1691 36 1693 38
rect 1786 44 1788 46
rect 1705 36 1707 38
rect 1826 44 1828 46
rect 1796 37 1798 39
rect 1866 49 1868 51
rect 1836 36 1838 38
rect 1931 44 1933 46
rect 1850 36 1852 38
rect 1971 49 1973 51
rect 1941 36 1943 38
rect 1955 36 1957 38
<< ndifct0 >>
rect 35 214 37 216
rect 75 214 77 216
rect 150 212 152 214
rect 162 215 164 217
rect 187 214 189 216
rect 176 207 178 209
rect 395 213 397 215
rect 405 213 407 215
rect 475 213 477 215
rect 500 214 502 216
rect 486 206 488 208
rect 512 211 514 213
rect 600 213 602 215
rect 610 213 612 215
rect 680 213 682 215
rect 705 214 707 216
rect 691 206 693 208
rect 717 211 719 213
rect 1825 214 1827 216
rect 1865 214 1867 216
rect 1940 212 1942 214
rect 1952 215 1954 217
rect 1977 214 1979 216
rect 1966 207 1968 209
rect 65 102 67 104
rect 75 102 77 104
rect 156 109 158 111
rect 145 102 147 104
rect 170 101 172 103
rect 182 104 184 106
rect 280 109 282 111
rect 269 102 271 104
rect 294 101 296 103
rect 306 104 308 106
rect 365 101 367 103
rect 405 101 407 103
rect 480 103 482 105
rect 506 108 508 110
rect 492 100 494 102
rect 517 101 519 103
rect 570 101 572 103
rect 610 101 612 103
rect 685 103 687 105
rect 711 108 713 110
rect 697 100 699 102
rect 722 101 724 103
rect 797 109 799 111
rect 788 96 790 98
rect 858 109 860 111
rect 847 102 849 104
rect 872 101 874 103
rect 807 96 809 98
rect 884 104 886 106
rect 963 109 965 111
rect 952 102 954 104
rect 977 101 979 103
rect 989 104 991 106
rect 1047 109 1049 111
rect 1038 96 1040 98
rect 1108 109 1110 111
rect 1097 102 1099 104
rect 1122 101 1124 103
rect 1057 96 1059 98
rect 1134 104 1136 106
rect 1213 109 1215 111
rect 1202 102 1204 104
rect 1227 101 1229 103
rect 1239 104 1241 106
rect 1297 109 1299 111
rect 1288 96 1290 98
rect 1358 109 1360 111
rect 1347 102 1349 104
rect 1372 101 1374 103
rect 1307 96 1309 98
rect 1384 104 1386 106
rect 1463 109 1465 111
rect 1452 102 1454 104
rect 1477 101 1479 103
rect 1489 104 1491 106
rect 1547 109 1549 111
rect 1538 96 1540 98
rect 1608 109 1610 111
rect 1597 102 1599 104
rect 1622 101 1624 103
rect 1557 96 1559 98
rect 1634 104 1636 106
rect 1713 109 1715 111
rect 1702 102 1704 104
rect 1727 101 1729 103
rect 1739 104 1741 106
rect 1855 102 1857 104
rect 1865 102 1867 104
rect 1946 109 1948 111
rect 1935 102 1937 104
rect 1960 101 1962 103
rect 1972 104 1974 106
rect 20 66 22 68
rect 39 66 41 68
rect 29 53 31 55
rect 79 60 81 62
rect 104 61 106 63
rect 90 53 92 55
rect 116 58 118 60
rect 184 60 186 62
rect 209 61 211 63
rect 195 53 197 55
rect 221 58 223 60
rect 270 66 272 68
rect 289 66 291 68
rect 279 53 281 55
rect 329 60 331 62
rect 354 61 356 63
rect 340 53 342 55
rect 366 58 368 60
rect 434 60 436 62
rect 459 61 461 63
rect 445 53 447 55
rect 471 58 473 60
rect 520 66 522 68
rect 539 66 541 68
rect 529 53 531 55
rect 579 60 581 62
rect 604 61 606 63
rect 590 53 592 55
rect 616 58 618 60
rect 684 60 686 62
rect 709 61 711 63
rect 695 53 697 55
rect 721 58 723 60
rect 770 66 772 68
rect 789 66 791 68
rect 779 53 781 55
rect 829 60 831 62
rect 854 61 856 63
rect 840 53 842 55
rect 866 58 868 60
rect 934 60 936 62
rect 959 61 961 63
rect 945 53 947 55
rect 971 58 973 60
rect 1030 66 1032 68
rect 1049 66 1051 68
rect 1039 53 1041 55
rect 1089 60 1091 62
rect 1114 61 1116 63
rect 1100 53 1102 55
rect 1126 58 1128 60
rect 1194 60 1196 62
rect 1219 61 1221 63
rect 1205 53 1207 55
rect 1231 58 1233 60
rect 1280 66 1282 68
rect 1299 66 1301 68
rect 1289 53 1291 55
rect 1339 60 1341 62
rect 1364 61 1366 63
rect 1350 53 1352 55
rect 1376 58 1378 60
rect 1444 60 1446 62
rect 1469 61 1471 63
rect 1455 53 1457 55
rect 1481 58 1483 60
rect 1530 66 1532 68
rect 1549 66 1551 68
rect 1539 53 1541 55
rect 1589 60 1591 62
rect 1614 61 1616 63
rect 1600 53 1602 55
rect 1626 58 1628 60
rect 1694 60 1696 62
rect 1719 61 1721 63
rect 1705 53 1707 55
rect 1731 58 1733 60
rect 1780 66 1782 68
rect 1799 66 1801 68
rect 1789 53 1791 55
rect 1839 60 1841 62
rect 1864 61 1866 63
rect 1850 53 1852 55
rect 1876 58 1878 60
rect 1944 60 1946 62
rect 1969 61 1971 63
rect 1955 53 1957 55
rect 1981 58 1983 60
<< ndifct1 >>
rect 54 224 56 226
rect 94 224 96 226
rect 122 224 124 226
rect 65 212 67 214
rect 105 212 107 214
rect 206 224 208 226
rect 140 214 142 216
rect 376 223 378 225
rect 424 223 426 225
rect 456 223 458 225
rect 217 212 219 214
rect 365 211 367 213
rect 540 223 542 225
rect 581 223 583 225
rect 435 211 437 213
rect 445 211 447 213
rect 522 213 524 215
rect 629 223 631 225
rect 661 223 663 225
rect 570 211 572 213
rect 745 223 747 225
rect 1844 224 1846 226
rect 640 211 642 213
rect 650 211 652 213
rect 727 213 729 215
rect 1884 224 1886 226
rect 1912 224 1914 226
rect 1855 212 1857 214
rect 1895 212 1897 214
rect 1996 224 1998 226
rect 1930 214 1932 216
rect 2007 212 2009 214
rect 35 104 37 106
rect 105 104 107 106
rect 115 104 117 106
rect 46 92 48 94
rect 94 92 96 94
rect 192 102 194 104
rect 126 92 128 94
rect 239 104 241 106
rect 210 92 212 94
rect 316 102 318 104
rect 250 92 252 94
rect 395 103 397 105
rect 334 92 336 94
rect 435 103 437 105
rect 384 91 386 93
rect 470 101 472 103
rect 547 103 549 105
rect 424 91 426 93
rect 452 91 454 93
rect 600 103 602 105
rect 536 91 538 93
rect 640 103 642 105
rect 589 91 591 93
rect 675 101 677 103
rect 777 109 779 111
rect 752 103 754 105
rect 629 91 631 93
rect 657 91 659 93
rect 817 104 819 106
rect 741 91 743 93
rect 894 102 896 104
rect 828 92 830 94
rect 922 104 924 106
rect 1027 109 1029 111
rect 912 92 914 94
rect 999 102 1001 104
rect 933 92 935 94
rect 1067 104 1069 106
rect 1017 92 1019 94
rect 1144 102 1146 104
rect 1078 92 1080 94
rect 1172 104 1174 106
rect 1277 109 1279 111
rect 1162 92 1164 94
rect 1249 102 1251 104
rect 1183 92 1185 94
rect 1317 104 1319 106
rect 1267 92 1269 94
rect 1394 102 1396 104
rect 1328 92 1330 94
rect 1422 104 1424 106
rect 1527 109 1529 111
rect 1412 92 1414 94
rect 1499 102 1501 104
rect 1433 92 1435 94
rect 1567 104 1569 106
rect 1517 92 1519 94
rect 1644 102 1646 104
rect 1578 92 1580 94
rect 1672 104 1674 106
rect 1662 92 1664 94
rect 1749 102 1751 104
rect 1683 92 1685 94
rect 1825 104 1827 106
rect 1895 104 1897 106
rect 1905 104 1907 106
rect 1767 92 1769 94
rect 1836 92 1838 94
rect 1884 92 1886 94
rect 1982 102 1984 104
rect 1916 92 1918 94
rect 2000 92 2002 94
rect 60 70 62 72
rect 9 53 11 55
rect 144 70 146 72
rect 165 70 167 72
rect 49 58 51 60
rect 126 60 128 62
rect 249 70 251 72
rect 154 58 156 60
rect 231 60 233 62
rect 310 70 312 72
rect 259 53 261 55
rect 394 70 396 72
rect 415 70 417 72
rect 299 58 301 60
rect 376 60 378 62
rect 499 70 501 72
rect 404 58 406 60
rect 481 60 483 62
rect 560 70 562 72
rect 509 53 511 55
rect 644 70 646 72
rect 665 70 667 72
rect 549 58 551 60
rect 626 60 628 62
rect 749 70 751 72
rect 654 58 656 60
rect 731 60 733 62
rect 810 70 812 72
rect 759 53 761 55
rect 894 70 896 72
rect 915 70 917 72
rect 799 58 801 60
rect 876 60 878 62
rect 999 70 1001 72
rect 904 58 906 60
rect 981 60 983 62
rect 1070 70 1072 72
rect 1019 53 1021 55
rect 1154 70 1156 72
rect 1175 70 1177 72
rect 1059 58 1061 60
rect 1136 60 1138 62
rect 1259 70 1261 72
rect 1164 58 1166 60
rect 1241 60 1243 62
rect 1320 70 1322 72
rect 1269 53 1271 55
rect 1404 70 1406 72
rect 1425 70 1427 72
rect 1309 58 1311 60
rect 1386 60 1388 62
rect 1509 70 1511 72
rect 1414 58 1416 60
rect 1491 60 1493 62
rect 1570 70 1572 72
rect 1519 53 1521 55
rect 1654 70 1656 72
rect 1675 70 1677 72
rect 1559 58 1561 60
rect 1636 60 1638 62
rect 1759 70 1761 72
rect 1664 58 1666 60
rect 1741 60 1743 62
rect 1820 70 1822 72
rect 1769 53 1771 55
rect 1904 70 1906 72
rect 1925 70 1927 72
rect 1809 58 1811 60
rect 1886 60 1888 62
rect 2009 70 2011 72
rect 1914 58 1916 60
rect 1991 60 1993 62
<< ntiect1 >>
rect 64 164 66 166
rect 104 164 106 166
rect 142 164 144 166
rect 216 164 218 166
rect 366 163 368 165
rect 434 163 436 165
rect 446 163 448 165
rect 520 163 522 165
rect 571 163 573 165
rect 639 163 641 165
rect 651 163 653 165
rect 725 163 727 165
rect 1854 164 1856 166
rect 1894 164 1896 166
rect 1932 164 1934 166
rect 2006 164 2008 166
rect 36 152 38 154
rect 104 152 106 154
rect 116 152 118 154
rect 190 152 192 154
rect 240 152 242 154
rect 314 152 316 154
rect 394 151 396 153
rect 434 151 436 153
rect 472 151 474 153
rect 546 151 548 153
rect 599 151 601 153
rect 639 151 641 153
rect 677 151 679 153
rect 751 151 753 153
rect 778 152 780 154
rect 818 152 820 154
rect 892 152 894 154
rect 923 152 925 154
rect 997 152 999 154
rect 1028 152 1030 154
rect 1068 152 1070 154
rect 1142 152 1144 154
rect 1173 152 1175 154
rect 1247 152 1249 154
rect 1278 152 1280 154
rect 1318 152 1320 154
rect 1392 152 1394 154
rect 1423 152 1425 154
rect 1497 152 1499 154
rect 1528 152 1530 154
rect 1568 152 1570 154
rect 1642 152 1644 154
rect 1673 152 1675 154
rect 1747 152 1749 154
rect 1826 152 1828 154
rect 1894 152 1896 154
rect 1906 152 1908 154
rect 1980 152 1982 154
rect 10 10 12 12
rect 50 10 52 12
rect 124 10 126 12
rect 155 10 157 12
rect 229 10 231 12
rect 260 10 262 12
rect 300 10 302 12
rect 374 10 376 12
rect 405 10 407 12
rect 479 10 481 12
rect 510 10 512 12
rect 550 10 552 12
rect 624 10 626 12
rect 655 10 657 12
rect 729 10 731 12
rect 760 10 762 12
rect 800 10 802 12
rect 874 10 876 12
rect 905 10 907 12
rect 979 10 981 12
rect 1020 10 1022 12
rect 1060 10 1062 12
rect 1134 10 1136 12
rect 1165 10 1167 12
rect 1239 10 1241 12
rect 1270 10 1272 12
rect 1310 10 1312 12
rect 1384 10 1386 12
rect 1415 10 1417 12
rect 1489 10 1491 12
rect 1520 10 1522 12
rect 1560 10 1562 12
rect 1634 10 1636 12
rect 1665 10 1667 12
rect 1739 10 1741 12
rect 1770 10 1772 12
rect 1810 10 1812 12
rect 1884 10 1886 12
rect 1915 10 1917 12
rect 1989 10 1991 12
<< ptiect1 >>
rect 64 224 66 226
rect 104 224 106 226
rect 175 224 177 226
rect 216 224 218 226
rect 366 223 368 225
rect 434 223 436 225
rect 446 223 448 225
rect 487 223 489 225
rect 571 223 573 225
rect 639 223 641 225
rect 651 223 653 225
rect 692 223 694 225
rect 1854 224 1856 226
rect 1894 224 1896 226
rect 1965 224 1967 226
rect 2006 224 2008 226
rect 36 92 38 94
rect 104 92 106 94
rect 116 92 118 94
rect 157 92 159 94
rect 240 92 242 94
rect 281 92 283 94
rect 394 91 396 93
rect 434 91 436 93
rect 505 91 507 93
rect 546 91 548 93
rect 599 91 601 93
rect 639 91 641 93
rect 710 91 712 93
rect 751 91 753 93
rect 778 92 780 94
rect 818 92 820 94
rect 859 92 861 94
rect 923 92 925 94
rect 964 92 966 94
rect 1028 92 1030 94
rect 1068 92 1070 94
rect 1109 92 1111 94
rect 1173 92 1175 94
rect 1214 92 1216 94
rect 1278 92 1280 94
rect 1318 92 1320 94
rect 1359 92 1361 94
rect 1423 92 1425 94
rect 1464 92 1466 94
rect 1528 92 1530 94
rect 1568 92 1570 94
rect 1609 92 1611 94
rect 1673 92 1675 94
rect 1714 92 1716 94
rect 1826 92 1828 94
rect 1894 92 1896 94
rect 1906 92 1908 94
rect 1947 92 1949 94
rect 10 70 12 72
rect 50 70 52 72
rect 91 70 93 72
rect 155 70 157 72
rect 196 70 198 72
rect 260 70 262 72
rect 300 70 302 72
rect 341 70 343 72
rect 405 70 407 72
rect 446 70 448 72
rect 510 70 512 72
rect 550 70 552 72
rect 591 70 593 72
rect 655 70 657 72
rect 696 70 698 72
rect 760 70 762 72
rect 800 70 802 72
rect 841 70 843 72
rect 905 70 907 72
rect 946 70 948 72
rect 1020 70 1022 72
rect 1060 70 1062 72
rect 1101 70 1103 72
rect 1165 70 1167 72
rect 1206 70 1208 72
rect 1270 70 1272 72
rect 1310 70 1312 72
rect 1351 70 1353 72
rect 1415 70 1417 72
rect 1456 70 1458 72
rect 1520 70 1522 72
rect 1560 70 1562 72
rect 1601 70 1603 72
rect 1665 70 1667 72
rect 1706 70 1708 72
rect 1770 70 1772 72
rect 1810 70 1812 72
rect 1851 70 1853 72
rect 1915 70 1917 72
rect 1956 70 1958 72
<< pdifct0 >>
rect 35 174 37 176
rect 45 181 47 183
rect 45 174 47 176
rect 55 176 57 178
rect 75 174 77 176
rect 85 181 87 183
rect 85 174 87 176
rect 95 176 97 178
rect 122 173 124 175
rect 142 188 144 190
rect 142 181 144 183
rect 158 174 160 176
rect 158 167 160 169
rect 168 188 170 190
rect 187 174 189 176
rect 197 181 199 183
rect 197 174 199 176
rect 207 176 209 178
rect 375 175 377 177
rect 385 180 387 182
rect 385 173 387 175
rect 395 173 397 175
rect 405 173 407 175
rect 415 180 417 182
rect 415 173 417 175
rect 425 175 427 177
rect 494 187 496 189
rect 455 175 457 177
rect 465 180 467 182
rect 465 173 467 175
rect 475 173 477 175
rect 504 173 506 175
rect 520 187 522 189
rect 520 180 522 182
rect 504 166 506 168
rect 540 172 542 174
rect 580 175 582 177
rect 590 180 592 182
rect 590 173 592 175
rect 600 173 602 175
rect 610 173 612 175
rect 620 180 622 182
rect 620 173 622 175
rect 630 175 632 177
rect 699 187 701 189
rect 660 175 662 177
rect 670 180 672 182
rect 670 173 672 175
rect 680 173 682 175
rect 709 173 711 175
rect 725 187 727 189
rect 725 180 727 182
rect 709 166 711 168
rect 745 172 747 174
rect 1825 174 1827 176
rect 1835 181 1837 183
rect 1835 174 1837 176
rect 1845 176 1847 178
rect 1865 174 1867 176
rect 1875 181 1877 183
rect 1875 174 1877 176
rect 1885 176 1887 178
rect 1912 173 1914 175
rect 1932 188 1934 190
rect 1932 181 1934 183
rect 1948 174 1950 176
rect 1948 167 1950 169
rect 1958 188 1960 190
rect 1977 174 1979 176
rect 1987 181 1989 183
rect 1987 174 1989 176
rect 1997 176 1999 178
rect 45 140 47 142
rect 55 142 57 144
rect 55 135 57 137
rect 65 142 67 144
rect 75 142 77 144
rect 85 142 87 144
rect 85 135 87 137
rect 95 140 97 142
rect 125 140 127 142
rect 135 142 137 144
rect 135 135 137 137
rect 145 142 147 144
rect 164 128 166 130
rect 174 149 176 151
rect 174 142 176 144
rect 190 135 192 137
rect 190 128 192 130
rect 210 143 212 145
rect 249 140 251 142
rect 259 142 261 144
rect 259 135 261 137
rect 269 142 271 144
rect 288 128 290 130
rect 298 149 300 151
rect 298 142 300 144
rect 314 135 316 137
rect 314 128 316 130
rect 334 143 336 145
rect 365 141 367 143
rect 375 141 377 143
rect 375 134 377 136
rect 385 139 387 141
rect 405 141 407 143
rect 415 141 417 143
rect 415 134 417 136
rect 425 139 427 141
rect 452 142 454 144
rect 488 148 490 150
rect 472 134 474 136
rect 472 127 474 129
rect 488 141 490 143
rect 517 141 519 143
rect 527 141 529 143
rect 527 134 529 136
rect 537 139 539 141
rect 498 127 500 129
rect 570 141 572 143
rect 580 141 582 143
rect 580 134 582 136
rect 590 139 592 141
rect 610 141 612 143
rect 620 141 622 143
rect 620 134 622 136
rect 630 139 632 141
rect 657 142 659 144
rect 693 148 695 150
rect 677 134 679 136
rect 677 127 679 129
rect 693 141 695 143
rect 788 149 790 151
rect 722 141 724 143
rect 732 141 734 143
rect 732 134 734 136
rect 742 139 744 141
rect 703 127 705 129
rect 807 142 809 144
rect 827 140 829 142
rect 837 142 839 144
rect 837 135 839 137
rect 847 142 849 144
rect 866 128 868 130
rect 876 149 878 151
rect 876 142 878 144
rect 892 135 894 137
rect 892 128 894 130
rect 912 143 914 145
rect 932 140 934 142
rect 942 142 944 144
rect 942 135 944 137
rect 952 142 954 144
rect 971 128 973 130
rect 981 149 983 151
rect 981 142 983 144
rect 997 135 999 137
rect 997 128 999 130
rect 1038 149 1040 151
rect 1017 143 1019 145
rect 1057 142 1059 144
rect 1077 140 1079 142
rect 1087 142 1089 144
rect 1087 135 1089 137
rect 1097 142 1099 144
rect 1116 128 1118 130
rect 1126 149 1128 151
rect 1126 142 1128 144
rect 1142 135 1144 137
rect 1142 128 1144 130
rect 1162 143 1164 145
rect 1182 140 1184 142
rect 1192 142 1194 144
rect 1192 135 1194 137
rect 1202 142 1204 144
rect 1221 128 1223 130
rect 1231 149 1233 151
rect 1231 142 1233 144
rect 1247 135 1249 137
rect 1247 128 1249 130
rect 1288 149 1290 151
rect 1267 143 1269 145
rect 1307 142 1309 144
rect 1327 140 1329 142
rect 1337 142 1339 144
rect 1337 135 1339 137
rect 1347 142 1349 144
rect 1366 128 1368 130
rect 1376 149 1378 151
rect 1376 142 1378 144
rect 1392 135 1394 137
rect 1392 128 1394 130
rect 1412 143 1414 145
rect 1432 140 1434 142
rect 1442 142 1444 144
rect 1442 135 1444 137
rect 1452 142 1454 144
rect 1471 128 1473 130
rect 1481 149 1483 151
rect 1481 142 1483 144
rect 1497 135 1499 137
rect 1497 128 1499 130
rect 1538 149 1540 151
rect 1517 143 1519 145
rect 1557 142 1559 144
rect 1577 140 1579 142
rect 1587 142 1589 144
rect 1587 135 1589 137
rect 1597 142 1599 144
rect 1616 128 1618 130
rect 1626 149 1628 151
rect 1626 142 1628 144
rect 1642 135 1644 137
rect 1642 128 1644 130
rect 1662 143 1664 145
rect 1682 140 1684 142
rect 1692 142 1694 144
rect 1692 135 1694 137
rect 1702 142 1704 144
rect 1721 128 1723 130
rect 1731 149 1733 151
rect 1731 142 1733 144
rect 1747 135 1749 137
rect 1747 128 1749 130
rect 1767 143 1769 145
rect 1835 140 1837 142
rect 1845 142 1847 144
rect 1845 135 1847 137
rect 1855 142 1857 144
rect 1865 142 1867 144
rect 1875 142 1877 144
rect 1875 135 1877 137
rect 1885 140 1887 142
rect 1915 140 1917 142
rect 1925 142 1927 144
rect 1925 135 1927 137
rect 1935 142 1937 144
rect 1954 128 1956 130
rect 1964 149 1966 151
rect 1964 142 1966 144
rect 1980 135 1982 137
rect 1980 128 1982 130
rect 2000 143 2002 145
rect 20 13 22 15
rect 39 20 41 22
rect 98 34 100 36
rect 59 22 61 24
rect 69 27 71 29
rect 69 20 71 22
rect 79 20 81 22
rect 108 20 110 22
rect 124 34 126 36
rect 124 27 126 29
rect 108 13 110 15
rect 144 19 146 21
rect 203 34 205 36
rect 164 22 166 24
rect 174 27 176 29
rect 174 20 176 22
rect 184 20 186 22
rect 213 20 215 22
rect 229 34 231 36
rect 229 27 231 29
rect 213 13 215 15
rect 249 19 251 21
rect 270 13 272 15
rect 289 20 291 22
rect 348 34 350 36
rect 309 22 311 24
rect 319 27 321 29
rect 319 20 321 22
rect 329 20 331 22
rect 358 20 360 22
rect 374 34 376 36
rect 374 27 376 29
rect 358 13 360 15
rect 394 19 396 21
rect 453 34 455 36
rect 414 22 416 24
rect 424 27 426 29
rect 424 20 426 22
rect 434 20 436 22
rect 463 20 465 22
rect 479 34 481 36
rect 479 27 481 29
rect 463 13 465 15
rect 499 19 501 21
rect 520 13 522 15
rect 539 20 541 22
rect 598 34 600 36
rect 559 22 561 24
rect 569 27 571 29
rect 569 20 571 22
rect 579 20 581 22
rect 608 20 610 22
rect 624 34 626 36
rect 624 27 626 29
rect 608 13 610 15
rect 644 19 646 21
rect 703 34 705 36
rect 664 22 666 24
rect 674 27 676 29
rect 674 20 676 22
rect 684 20 686 22
rect 713 20 715 22
rect 729 34 731 36
rect 729 27 731 29
rect 713 13 715 15
rect 749 19 751 21
rect 770 13 772 15
rect 789 20 791 22
rect 848 34 850 36
rect 809 22 811 24
rect 819 27 821 29
rect 819 20 821 22
rect 829 20 831 22
rect 858 20 860 22
rect 874 34 876 36
rect 874 27 876 29
rect 858 13 860 15
rect 894 19 896 21
rect 953 34 955 36
rect 914 22 916 24
rect 924 27 926 29
rect 924 20 926 22
rect 934 20 936 22
rect 963 20 965 22
rect 979 34 981 36
rect 979 27 981 29
rect 963 13 965 15
rect 999 19 1001 21
rect 1030 13 1032 15
rect 1049 20 1051 22
rect 1108 34 1110 36
rect 1069 22 1071 24
rect 1079 27 1081 29
rect 1079 20 1081 22
rect 1089 20 1091 22
rect 1118 20 1120 22
rect 1134 34 1136 36
rect 1134 27 1136 29
rect 1118 13 1120 15
rect 1154 19 1156 21
rect 1213 34 1215 36
rect 1174 22 1176 24
rect 1184 27 1186 29
rect 1184 20 1186 22
rect 1194 20 1196 22
rect 1223 20 1225 22
rect 1239 34 1241 36
rect 1239 27 1241 29
rect 1223 13 1225 15
rect 1259 19 1261 21
rect 1280 13 1282 15
rect 1299 20 1301 22
rect 1358 34 1360 36
rect 1319 22 1321 24
rect 1329 27 1331 29
rect 1329 20 1331 22
rect 1339 20 1341 22
rect 1368 20 1370 22
rect 1384 34 1386 36
rect 1384 27 1386 29
rect 1368 13 1370 15
rect 1404 19 1406 21
rect 1463 34 1465 36
rect 1424 22 1426 24
rect 1434 27 1436 29
rect 1434 20 1436 22
rect 1444 20 1446 22
rect 1473 20 1475 22
rect 1489 34 1491 36
rect 1489 27 1491 29
rect 1473 13 1475 15
rect 1509 19 1511 21
rect 1530 13 1532 15
rect 1549 20 1551 22
rect 1608 34 1610 36
rect 1569 22 1571 24
rect 1579 27 1581 29
rect 1579 20 1581 22
rect 1589 20 1591 22
rect 1618 20 1620 22
rect 1634 34 1636 36
rect 1634 27 1636 29
rect 1618 13 1620 15
rect 1654 19 1656 21
rect 1713 34 1715 36
rect 1674 22 1676 24
rect 1684 27 1686 29
rect 1684 20 1686 22
rect 1694 20 1696 22
rect 1723 20 1725 22
rect 1739 34 1741 36
rect 1739 27 1741 29
rect 1723 13 1725 15
rect 1759 19 1761 21
rect 1780 13 1782 15
rect 1799 20 1801 22
rect 1858 34 1860 36
rect 1819 22 1821 24
rect 1829 27 1831 29
rect 1829 20 1831 22
rect 1839 20 1841 22
rect 1868 20 1870 22
rect 1884 34 1886 36
rect 1884 27 1886 29
rect 1868 13 1870 15
rect 1904 19 1906 21
rect 1963 34 1965 36
rect 1924 22 1926 24
rect 1934 27 1936 29
rect 1934 20 1936 22
rect 1944 20 1946 22
rect 1973 20 1975 22
rect 1989 34 1991 36
rect 1989 27 1991 29
rect 1973 13 1975 15
rect 2009 19 2011 21
<< pdifct1 >>
rect 65 188 67 190
rect 65 181 67 183
rect 105 188 107 190
rect 105 181 107 183
rect 132 181 134 183
rect 217 188 219 190
rect 217 181 219 183
rect 365 187 367 189
rect 365 180 367 182
rect 435 187 437 189
rect 435 180 437 182
rect 445 187 447 189
rect 445 180 447 182
rect 530 180 532 182
rect 570 187 572 189
rect 570 180 572 182
rect 640 187 642 189
rect 640 180 642 182
rect 650 187 652 189
rect 650 180 652 182
rect 735 180 737 182
rect 1855 188 1857 190
rect 1855 181 1857 183
rect 1895 188 1897 190
rect 1895 181 1897 183
rect 1922 181 1924 183
rect 2007 188 2009 190
rect 2007 181 2009 183
rect 35 135 37 137
rect 35 128 37 130
rect 105 135 107 137
rect 105 128 107 130
rect 115 135 117 137
rect 115 128 117 130
rect 200 135 202 137
rect 239 135 241 137
rect 239 128 241 130
rect 324 135 326 137
rect 395 134 397 136
rect 395 127 397 129
rect 435 134 437 136
rect 435 127 437 129
rect 462 134 464 136
rect 547 134 549 136
rect 547 127 549 129
rect 600 134 602 136
rect 600 127 602 129
rect 640 134 642 136
rect 640 127 642 129
rect 667 134 669 136
rect 777 139 779 141
rect 752 134 754 136
rect 777 132 779 134
rect 752 127 754 129
rect 817 135 819 137
rect 817 128 819 130
rect 902 135 904 137
rect 922 135 924 137
rect 922 128 924 130
rect 1007 135 1009 137
rect 1027 139 1029 141
rect 1027 132 1029 134
rect 1067 135 1069 137
rect 1067 128 1069 130
rect 1152 135 1154 137
rect 1172 135 1174 137
rect 1172 128 1174 130
rect 1257 135 1259 137
rect 1277 139 1279 141
rect 1277 132 1279 134
rect 1317 135 1319 137
rect 1317 128 1319 130
rect 1402 135 1404 137
rect 1422 135 1424 137
rect 1422 128 1424 130
rect 1507 135 1509 137
rect 1527 139 1529 141
rect 1527 132 1529 134
rect 1567 135 1569 137
rect 1567 128 1569 130
rect 1652 135 1654 137
rect 1672 135 1674 137
rect 1672 128 1674 130
rect 1757 135 1759 137
rect 1825 135 1827 137
rect 1825 128 1827 130
rect 1895 135 1897 137
rect 1895 128 1897 130
rect 1905 135 1907 137
rect 1905 128 1907 130
rect 1990 135 1992 137
rect 9 30 11 32
rect 9 23 11 25
rect 49 34 51 36
rect 49 27 51 29
rect 134 27 136 29
rect 154 34 156 36
rect 154 27 156 29
rect 239 27 241 29
rect 259 30 261 32
rect 259 23 261 25
rect 299 34 301 36
rect 299 27 301 29
rect 384 27 386 29
rect 404 34 406 36
rect 404 27 406 29
rect 489 27 491 29
rect 509 30 511 32
rect 509 23 511 25
rect 549 34 551 36
rect 549 27 551 29
rect 634 27 636 29
rect 654 34 656 36
rect 654 27 656 29
rect 739 27 741 29
rect 759 30 761 32
rect 759 23 761 25
rect 799 34 801 36
rect 799 27 801 29
rect 884 27 886 29
rect 904 34 906 36
rect 904 27 906 29
rect 989 27 991 29
rect 1019 30 1021 32
rect 1019 23 1021 25
rect 1059 34 1061 36
rect 1059 27 1061 29
rect 1144 27 1146 29
rect 1164 34 1166 36
rect 1164 27 1166 29
rect 1249 27 1251 29
rect 1269 30 1271 32
rect 1269 23 1271 25
rect 1309 34 1311 36
rect 1309 27 1311 29
rect 1394 27 1396 29
rect 1414 34 1416 36
rect 1414 27 1416 29
rect 1499 27 1501 29
rect 1519 30 1521 32
rect 1519 23 1521 25
rect 1559 34 1561 36
rect 1559 27 1561 29
rect 1644 27 1646 29
rect 1664 34 1666 36
rect 1664 27 1666 29
rect 1749 27 1751 29
rect 1769 30 1771 32
rect 1769 23 1771 25
rect 1809 34 1811 36
rect 1809 27 1811 29
rect 1894 27 1896 29
rect 1914 34 1916 36
rect 1914 27 1916 29
rect 1999 27 2001 29
<< alu0 >>
rect 33 216 53 217
rect 33 214 35 216
rect 37 214 53 216
rect 33 213 53 214
rect 49 209 53 213
rect 73 216 93 217
rect 73 214 75 216
rect 77 214 93 216
rect 73 213 93 214
rect 64 210 65 212
rect 49 205 61 209
rect 57 200 61 205
rect 57 198 58 200
rect 60 198 61 200
rect 57 186 61 198
rect 89 209 93 213
rect 160 217 166 223
rect 104 210 105 212
rect 89 205 101 209
rect 97 200 101 205
rect 97 198 98 200
rect 100 198 101 200
rect 44 183 61 186
rect 44 181 45 183
rect 47 182 61 183
rect 47 181 48 182
rect 33 176 39 177
rect 33 174 35 176
rect 37 174 39 176
rect 33 167 39 174
rect 44 176 48 181
rect 97 186 101 198
rect 84 183 101 186
rect 84 181 85 183
rect 87 182 101 183
rect 87 181 88 182
rect 44 174 45 176
rect 47 174 48 176
rect 44 172 48 174
rect 53 178 59 179
rect 53 176 55 178
rect 57 176 59 178
rect 53 167 59 176
rect 73 176 79 177
rect 73 174 75 176
rect 77 174 79 176
rect 73 167 79 174
rect 84 176 88 181
rect 149 214 153 216
rect 160 215 162 217
rect 164 215 166 217
rect 160 214 166 215
rect 185 216 205 217
rect 185 214 187 216
rect 189 214 205 216
rect 149 212 150 214
rect 152 212 153 214
rect 185 213 205 214
rect 149 209 153 212
rect 129 205 153 209
rect 129 201 133 205
rect 175 209 179 211
rect 175 207 176 209
rect 178 207 179 209
rect 128 199 133 201
rect 128 197 129 199
rect 131 197 133 199
rect 137 200 153 201
rect 137 198 139 200
rect 141 198 153 200
rect 137 197 153 198
rect 128 195 133 197
rect 129 193 133 195
rect 129 190 145 193
rect 129 189 142 190
rect 141 188 142 189
rect 144 188 145 190
rect 141 183 145 188
rect 141 181 142 183
rect 144 181 145 183
rect 141 179 145 181
rect 149 191 153 197
rect 175 201 179 207
rect 168 197 179 201
rect 201 209 205 213
rect 216 210 217 212
rect 201 205 213 209
rect 209 200 213 205
rect 209 198 210 200
rect 212 198 213 200
rect 168 191 172 197
rect 149 190 172 191
rect 149 188 168 190
rect 170 188 172 190
rect 149 187 172 188
rect 84 174 85 176
rect 87 174 88 176
rect 84 172 88 174
rect 93 178 99 179
rect 93 176 95 178
rect 97 176 99 178
rect 149 176 153 187
rect 209 186 213 198
rect 196 183 213 186
rect 196 181 197 183
rect 199 182 213 183
rect 199 181 200 182
rect 93 167 99 176
rect 120 175 153 176
rect 120 173 122 175
rect 124 173 153 175
rect 120 172 153 173
rect 157 176 161 178
rect 157 174 158 176
rect 160 174 161 176
rect 157 169 161 174
rect 185 176 191 177
rect 185 174 187 176
rect 189 174 191 176
rect 157 167 158 169
rect 160 167 161 169
rect 185 167 191 174
rect 196 176 200 181
rect 379 215 399 216
rect 379 213 395 215
rect 397 213 399 215
rect 379 212 399 213
rect 403 215 423 216
rect 403 213 405 215
rect 407 213 423 215
rect 403 212 423 213
rect 367 209 368 211
rect 379 208 383 212
rect 371 204 383 208
rect 371 199 375 204
rect 371 197 372 199
rect 374 197 375 199
rect 371 185 375 197
rect 419 208 423 212
rect 434 209 435 211
rect 419 204 431 208
rect 427 199 431 204
rect 427 197 428 199
rect 430 197 431 199
rect 371 182 388 185
rect 371 181 385 182
rect 196 174 197 176
rect 199 174 200 176
rect 196 172 200 174
rect 205 178 211 179
rect 384 180 385 181
rect 387 180 388 182
rect 205 176 207 178
rect 209 176 211 178
rect 205 167 211 176
rect 373 177 379 178
rect 373 175 375 177
rect 377 175 379 177
rect 373 166 379 175
rect 384 175 388 180
rect 427 185 431 197
rect 414 182 431 185
rect 414 180 415 182
rect 417 181 431 182
rect 417 180 418 181
rect 384 173 385 175
rect 387 173 388 175
rect 384 171 388 173
rect 393 175 399 176
rect 393 173 395 175
rect 397 173 399 175
rect 393 166 399 173
rect 403 175 409 176
rect 403 173 405 175
rect 407 173 409 175
rect 403 166 409 173
rect 414 175 418 180
rect 498 216 504 222
rect 459 215 479 216
rect 459 213 475 215
rect 477 213 479 215
rect 498 214 500 216
rect 502 214 504 216
rect 498 213 504 214
rect 511 213 515 215
rect 459 212 479 213
rect 447 209 448 211
rect 459 208 463 212
rect 511 211 512 213
rect 514 211 515 213
rect 451 204 463 208
rect 451 199 455 204
rect 451 197 452 199
rect 454 197 455 199
rect 451 185 455 197
rect 485 208 489 210
rect 485 206 486 208
rect 488 206 489 208
rect 485 200 489 206
rect 511 208 515 211
rect 511 204 535 208
rect 485 196 496 200
rect 492 190 496 196
rect 531 200 535 204
rect 511 199 527 200
rect 511 197 523 199
rect 525 197 527 199
rect 511 196 527 197
rect 531 198 536 200
rect 531 196 533 198
rect 535 196 536 198
rect 511 190 515 196
rect 531 194 536 196
rect 531 192 535 194
rect 492 189 515 190
rect 492 187 494 189
rect 496 187 515 189
rect 492 186 515 187
rect 451 182 468 185
rect 451 181 465 182
rect 464 180 465 181
rect 467 180 468 182
rect 414 173 415 175
rect 417 173 418 175
rect 414 171 418 173
rect 423 177 429 178
rect 423 175 425 177
rect 427 175 429 177
rect 423 166 429 175
rect 453 177 459 178
rect 453 175 455 177
rect 457 175 459 177
rect 453 166 459 175
rect 464 175 468 180
rect 464 173 465 175
rect 467 173 468 175
rect 464 171 468 173
rect 473 175 479 176
rect 473 173 475 175
rect 477 173 479 175
rect 473 166 479 173
rect 503 175 507 177
rect 503 173 504 175
rect 506 173 507 175
rect 503 168 507 173
rect 511 175 515 186
rect 519 189 535 192
rect 519 187 520 189
rect 522 188 535 189
rect 522 187 523 188
rect 519 182 523 187
rect 519 180 520 182
rect 522 180 523 182
rect 519 178 523 180
rect 584 215 604 216
rect 584 213 600 215
rect 602 213 604 215
rect 584 212 604 213
rect 608 215 628 216
rect 608 213 610 215
rect 612 213 628 215
rect 608 212 628 213
rect 572 209 573 211
rect 584 208 588 212
rect 576 204 588 208
rect 576 199 580 204
rect 576 197 577 199
rect 579 197 580 199
rect 576 185 580 197
rect 624 208 628 212
rect 639 209 640 211
rect 624 204 636 208
rect 632 199 636 204
rect 632 197 633 199
rect 635 197 636 199
rect 576 182 593 185
rect 576 181 590 182
rect 589 180 590 181
rect 592 180 593 182
rect 578 177 584 178
rect 578 175 580 177
rect 582 175 584 177
rect 511 174 544 175
rect 511 172 540 174
rect 542 172 544 174
rect 511 171 544 172
rect 503 166 504 168
rect 506 166 507 168
rect 578 166 584 175
rect 589 175 593 180
rect 632 185 636 197
rect 619 182 636 185
rect 619 180 620 182
rect 622 181 636 182
rect 622 180 623 181
rect 589 173 590 175
rect 592 173 593 175
rect 589 171 593 173
rect 598 175 604 176
rect 598 173 600 175
rect 602 173 604 175
rect 598 166 604 173
rect 608 175 614 176
rect 608 173 610 175
rect 612 173 614 175
rect 608 166 614 173
rect 619 175 623 180
rect 703 216 709 222
rect 1823 216 1843 217
rect 664 215 684 216
rect 664 213 680 215
rect 682 213 684 215
rect 703 214 705 216
rect 707 214 709 216
rect 703 213 709 214
rect 716 213 720 215
rect 664 212 684 213
rect 652 209 653 211
rect 664 208 668 212
rect 716 211 717 213
rect 719 211 720 213
rect 1823 214 1825 216
rect 1827 214 1843 216
rect 1823 213 1843 214
rect 656 204 668 208
rect 656 199 660 204
rect 656 197 657 199
rect 659 197 660 199
rect 656 185 660 197
rect 690 208 694 210
rect 690 206 691 208
rect 693 206 694 208
rect 690 200 694 206
rect 716 208 720 211
rect 716 204 740 208
rect 690 196 701 200
rect 697 190 701 196
rect 736 200 740 204
rect 716 199 732 200
rect 716 197 728 199
rect 730 197 732 199
rect 716 196 732 197
rect 736 198 741 200
rect 736 196 738 198
rect 740 196 741 198
rect 716 190 720 196
rect 736 194 741 196
rect 736 192 740 194
rect 697 189 720 190
rect 697 187 699 189
rect 701 187 720 189
rect 697 186 720 187
rect 656 182 673 185
rect 656 181 670 182
rect 669 180 670 181
rect 672 180 673 182
rect 619 173 620 175
rect 622 173 623 175
rect 619 171 623 173
rect 628 177 634 178
rect 628 175 630 177
rect 632 175 634 177
rect 628 166 634 175
rect 658 177 664 178
rect 658 175 660 177
rect 662 175 664 177
rect 658 166 664 175
rect 669 175 673 180
rect 669 173 670 175
rect 672 173 673 175
rect 669 171 673 173
rect 678 175 684 176
rect 678 173 680 175
rect 682 173 684 175
rect 678 166 684 173
rect 708 175 712 177
rect 708 173 709 175
rect 711 173 712 175
rect 708 168 712 173
rect 716 175 720 186
rect 724 189 740 192
rect 724 187 725 189
rect 727 188 740 189
rect 727 187 728 188
rect 724 182 728 187
rect 1839 209 1843 213
rect 1863 216 1883 217
rect 1863 214 1865 216
rect 1867 214 1883 216
rect 1863 213 1883 214
rect 1854 210 1855 212
rect 1839 205 1851 209
rect 1847 200 1851 205
rect 1847 198 1848 200
rect 1850 198 1851 200
rect 724 180 725 182
rect 727 180 728 182
rect 724 178 728 180
rect 1847 186 1851 198
rect 1879 209 1883 213
rect 1950 217 1956 223
rect 1894 210 1895 212
rect 1879 205 1891 209
rect 1887 200 1891 205
rect 1887 198 1888 200
rect 1890 198 1891 200
rect 1834 183 1851 186
rect 1834 181 1835 183
rect 1837 182 1851 183
rect 1837 181 1838 182
rect 1823 176 1829 177
rect 716 174 749 175
rect 716 172 745 174
rect 747 172 749 174
rect 716 171 749 172
rect 1823 174 1825 176
rect 1827 174 1829 176
rect 708 166 709 168
rect 711 166 712 168
rect 1823 167 1829 174
rect 1834 176 1838 181
rect 1887 186 1891 198
rect 1874 183 1891 186
rect 1874 181 1875 183
rect 1877 182 1891 183
rect 1877 181 1878 182
rect 1834 174 1835 176
rect 1837 174 1838 176
rect 1834 172 1838 174
rect 1843 178 1849 179
rect 1843 176 1845 178
rect 1847 176 1849 178
rect 1843 167 1849 176
rect 1863 176 1869 177
rect 1863 174 1865 176
rect 1867 174 1869 176
rect 1863 167 1869 174
rect 1874 176 1878 181
rect 1939 214 1943 216
rect 1950 215 1952 217
rect 1954 215 1956 217
rect 1950 214 1956 215
rect 1975 216 1995 217
rect 1975 214 1977 216
rect 1979 214 1995 216
rect 1939 212 1940 214
rect 1942 212 1943 214
rect 1975 213 1995 214
rect 1939 209 1943 212
rect 1919 205 1943 209
rect 1919 201 1923 205
rect 1965 209 1969 211
rect 1965 207 1966 209
rect 1968 207 1969 209
rect 1918 199 1923 201
rect 1918 197 1919 199
rect 1921 197 1923 199
rect 1927 200 1943 201
rect 1927 198 1929 200
rect 1931 198 1943 200
rect 1927 197 1943 198
rect 1918 195 1923 197
rect 1919 193 1923 195
rect 1919 190 1935 193
rect 1919 189 1932 190
rect 1931 188 1932 189
rect 1934 188 1935 190
rect 1931 183 1935 188
rect 1931 181 1932 183
rect 1934 181 1935 183
rect 1931 179 1935 181
rect 1939 191 1943 197
rect 1965 201 1969 207
rect 1958 197 1969 201
rect 1991 209 1995 213
rect 2006 210 2007 212
rect 1991 205 2003 209
rect 1999 200 2003 205
rect 1999 198 2000 200
rect 2002 198 2003 200
rect 1958 191 1962 197
rect 1939 190 1962 191
rect 1939 188 1958 190
rect 1960 188 1962 190
rect 1939 187 1962 188
rect 1874 174 1875 176
rect 1877 174 1878 176
rect 1874 172 1878 174
rect 1883 178 1889 179
rect 1883 176 1885 178
rect 1887 176 1889 178
rect 1939 176 1943 187
rect 1999 186 2003 198
rect 1986 183 2003 186
rect 1986 181 1987 183
rect 1989 182 2003 183
rect 1989 181 1990 182
rect 1883 167 1889 176
rect 1910 175 1943 176
rect 1910 173 1912 175
rect 1914 173 1943 175
rect 1910 172 1943 173
rect 1947 176 1951 178
rect 1947 174 1948 176
rect 1950 174 1951 176
rect 1947 169 1951 174
rect 1975 176 1981 177
rect 1975 174 1977 176
rect 1979 174 1981 176
rect 1947 167 1948 169
rect 1950 167 1951 169
rect 1975 167 1981 174
rect 1986 176 1990 181
rect 1986 174 1987 176
rect 1989 174 1990 176
rect 1986 172 1990 174
rect 1995 178 2001 179
rect 1995 176 1997 178
rect 1999 176 2001 178
rect 1995 167 2001 176
rect 43 142 49 151
rect 43 140 45 142
rect 47 140 49 142
rect 43 139 49 140
rect 54 144 58 146
rect 54 142 55 144
rect 57 142 58 144
rect 54 137 58 142
rect 63 144 69 151
rect 63 142 65 144
rect 67 142 69 144
rect 63 141 69 142
rect 73 144 79 151
rect 73 142 75 144
rect 77 142 79 144
rect 73 141 79 142
rect 84 144 88 146
rect 84 142 85 144
rect 87 142 88 144
rect 54 136 55 137
rect 41 135 55 136
rect 57 135 58 137
rect 41 132 58 135
rect 41 120 45 132
rect 84 137 88 142
rect 93 142 99 151
rect 93 140 95 142
rect 97 140 99 142
rect 93 139 99 140
rect 123 142 129 151
rect 123 140 125 142
rect 127 140 129 142
rect 123 139 129 140
rect 134 144 138 146
rect 134 142 135 144
rect 137 142 138 144
rect 84 135 85 137
rect 87 136 88 137
rect 87 135 101 136
rect 84 132 101 135
rect 41 118 42 120
rect 44 118 45 120
rect 41 113 45 118
rect 41 109 53 113
rect 37 106 38 108
rect 49 105 53 109
rect 97 120 101 132
rect 97 118 98 120
rect 100 118 101 120
rect 97 113 101 118
rect 89 109 101 113
rect 89 105 93 109
rect 104 106 105 108
rect 49 104 69 105
rect 49 102 65 104
rect 67 102 69 104
rect 49 101 69 102
rect 73 104 93 105
rect 73 102 75 104
rect 77 102 93 104
rect 73 101 93 102
rect 134 137 138 142
rect 143 144 149 151
rect 173 149 174 151
rect 176 149 177 151
rect 143 142 145 144
rect 147 142 149 144
rect 143 141 149 142
rect 173 144 177 149
rect 173 142 174 144
rect 176 142 177 144
rect 173 140 177 142
rect 181 145 214 146
rect 181 143 210 145
rect 212 143 214 145
rect 181 142 214 143
rect 247 142 253 151
rect 134 136 135 137
rect 121 135 135 136
rect 137 135 138 137
rect 121 132 138 135
rect 121 120 125 132
rect 181 131 185 142
rect 247 140 249 142
rect 251 140 253 142
rect 247 139 253 140
rect 258 144 262 146
rect 258 142 259 144
rect 261 142 262 144
rect 162 130 185 131
rect 162 128 164 130
rect 166 128 185 130
rect 162 127 185 128
rect 162 121 166 127
rect 121 118 122 120
rect 124 118 125 120
rect 121 113 125 118
rect 121 109 133 113
rect 117 106 118 108
rect 129 105 133 109
rect 155 117 166 121
rect 155 111 159 117
rect 181 121 185 127
rect 189 137 193 139
rect 189 135 190 137
rect 192 135 193 137
rect 189 130 193 135
rect 189 128 190 130
rect 192 129 193 130
rect 192 128 205 129
rect 189 125 205 128
rect 201 123 205 125
rect 201 121 206 123
rect 181 120 197 121
rect 181 118 193 120
rect 195 118 197 120
rect 181 117 197 118
rect 201 119 203 121
rect 205 119 206 121
rect 201 117 206 119
rect 155 109 156 111
rect 158 109 159 111
rect 155 107 159 109
rect 201 113 205 117
rect 181 109 205 113
rect 181 106 185 109
rect 129 104 149 105
rect 181 104 182 106
rect 184 104 185 106
rect 129 102 145 104
rect 147 102 149 104
rect 129 101 149 102
rect 168 103 174 104
rect 168 101 170 103
rect 172 101 174 103
rect 181 102 185 104
rect 258 137 262 142
rect 267 144 273 151
rect 297 149 298 151
rect 300 149 301 151
rect 267 142 269 144
rect 271 142 273 144
rect 267 141 273 142
rect 297 144 301 149
rect 297 142 298 144
rect 300 142 301 144
rect 297 140 301 142
rect 305 145 338 146
rect 305 143 334 145
rect 336 143 338 145
rect 305 142 338 143
rect 363 143 369 150
rect 258 136 259 137
rect 245 135 259 136
rect 261 135 262 137
rect 245 132 262 135
rect 245 120 249 132
rect 305 131 309 142
rect 363 141 365 143
rect 367 141 369 143
rect 363 140 369 141
rect 374 143 378 145
rect 374 141 375 143
rect 377 141 378 143
rect 286 130 309 131
rect 286 128 288 130
rect 290 128 309 130
rect 286 127 309 128
rect 286 121 290 127
rect 245 118 246 120
rect 248 118 249 120
rect 245 113 249 118
rect 245 109 257 113
rect 241 106 242 108
rect 168 95 174 101
rect 253 105 257 109
rect 279 117 290 121
rect 279 111 283 117
rect 305 121 309 127
rect 313 137 317 139
rect 313 135 314 137
rect 316 135 317 137
rect 313 130 317 135
rect 313 128 314 130
rect 316 129 317 130
rect 316 128 329 129
rect 313 125 329 128
rect 325 123 329 125
rect 325 121 330 123
rect 305 120 321 121
rect 305 118 317 120
rect 319 118 321 120
rect 305 117 321 118
rect 325 119 327 121
rect 329 119 330 121
rect 325 117 330 119
rect 279 109 280 111
rect 282 109 283 111
rect 279 107 283 109
rect 325 113 329 117
rect 305 109 329 113
rect 305 106 309 109
rect 253 104 273 105
rect 305 104 306 106
rect 308 104 309 106
rect 374 136 378 141
rect 383 141 389 150
rect 383 139 385 141
rect 387 139 389 141
rect 403 143 409 150
rect 403 141 405 143
rect 407 141 409 143
rect 403 140 409 141
rect 414 143 418 145
rect 414 141 415 143
rect 417 141 418 143
rect 383 138 389 139
rect 374 134 375 136
rect 377 135 378 136
rect 377 134 391 135
rect 374 131 391 134
rect 387 119 391 131
rect 387 117 388 119
rect 390 117 391 119
rect 387 112 391 117
rect 379 108 391 112
rect 414 136 418 141
rect 423 141 429 150
rect 487 148 488 150
rect 490 148 491 150
rect 450 144 483 145
rect 450 142 452 144
rect 454 142 483 144
rect 450 141 483 142
rect 423 139 425 141
rect 427 139 429 141
rect 423 138 429 139
rect 414 134 415 136
rect 417 135 418 136
rect 417 134 431 135
rect 414 131 431 134
rect 253 102 269 104
rect 271 102 273 104
rect 253 101 273 102
rect 292 103 298 104
rect 292 101 294 103
rect 296 101 298 103
rect 305 102 309 104
rect 379 104 383 108
rect 394 105 395 107
rect 427 119 431 131
rect 427 117 428 119
rect 430 117 431 119
rect 427 112 431 117
rect 419 108 431 112
rect 363 103 383 104
rect 363 101 365 103
rect 367 101 383 103
rect 292 95 298 101
rect 363 100 383 101
rect 419 104 423 108
rect 434 105 435 107
rect 403 103 423 104
rect 403 101 405 103
rect 407 101 423 103
rect 403 100 423 101
rect 471 136 475 138
rect 471 134 472 136
rect 474 134 475 136
rect 471 129 475 134
rect 471 128 472 129
rect 459 127 472 128
rect 474 127 475 129
rect 459 124 475 127
rect 479 130 483 141
rect 487 143 491 148
rect 487 141 488 143
rect 490 141 491 143
rect 487 139 491 141
rect 515 143 521 150
rect 515 141 517 143
rect 519 141 521 143
rect 515 140 521 141
rect 526 143 530 145
rect 526 141 527 143
rect 529 141 530 143
rect 526 136 530 141
rect 535 141 541 150
rect 535 139 537 141
rect 539 139 541 141
rect 568 143 574 150
rect 568 141 570 143
rect 572 141 574 143
rect 568 140 574 141
rect 579 143 583 145
rect 579 141 580 143
rect 582 141 583 143
rect 535 138 541 139
rect 526 134 527 136
rect 529 135 530 136
rect 529 134 543 135
rect 526 131 543 134
rect 479 129 502 130
rect 479 127 498 129
rect 500 127 502 129
rect 479 126 502 127
rect 459 122 463 124
rect 458 120 463 122
rect 479 120 483 126
rect 458 118 459 120
rect 461 118 463 120
rect 458 116 463 118
rect 467 119 483 120
rect 467 117 469 119
rect 471 117 483 119
rect 467 116 483 117
rect 459 112 463 116
rect 498 120 502 126
rect 498 116 509 120
rect 459 108 483 112
rect 479 105 483 108
rect 505 110 509 116
rect 505 108 506 110
rect 508 108 509 110
rect 505 106 509 108
rect 539 119 543 131
rect 539 117 540 119
rect 542 117 543 119
rect 539 112 543 117
rect 531 108 543 112
rect 579 136 583 141
rect 588 141 594 150
rect 588 139 590 141
rect 592 139 594 141
rect 608 143 614 150
rect 608 141 610 143
rect 612 141 614 143
rect 608 140 614 141
rect 619 143 623 145
rect 619 141 620 143
rect 622 141 623 143
rect 588 138 594 139
rect 579 134 580 136
rect 582 135 583 136
rect 582 134 596 135
rect 579 131 596 134
rect 479 103 480 105
rect 482 103 483 105
rect 531 104 535 108
rect 546 105 547 107
rect 592 119 596 131
rect 592 117 593 119
rect 595 117 596 119
rect 592 112 596 117
rect 584 108 596 112
rect 619 136 623 141
rect 628 141 634 150
rect 692 148 693 150
rect 695 148 696 150
rect 655 144 688 145
rect 655 142 657 144
rect 659 142 688 144
rect 655 141 688 142
rect 628 139 630 141
rect 632 139 634 141
rect 628 138 634 139
rect 619 134 620 136
rect 622 135 623 136
rect 622 134 636 135
rect 619 131 636 134
rect 515 103 535 104
rect 479 101 483 103
rect 490 102 496 103
rect 490 100 492 102
rect 494 100 496 102
rect 515 101 517 103
rect 519 101 535 103
rect 515 100 535 101
rect 584 104 588 108
rect 599 105 600 107
rect 632 119 636 131
rect 632 117 633 119
rect 635 117 636 119
rect 632 112 636 117
rect 624 108 636 112
rect 490 94 496 100
rect 568 103 588 104
rect 568 101 570 103
rect 572 101 588 103
rect 568 100 588 101
rect 624 104 628 108
rect 639 105 640 107
rect 608 103 628 104
rect 608 101 610 103
rect 612 101 628 103
rect 608 100 628 101
rect 676 136 680 138
rect 676 134 677 136
rect 679 134 680 136
rect 676 129 680 134
rect 676 128 677 129
rect 664 127 677 128
rect 679 127 680 129
rect 664 124 680 127
rect 684 130 688 141
rect 692 143 696 148
rect 692 141 693 143
rect 695 141 696 143
rect 692 139 696 141
rect 720 143 726 150
rect 720 141 722 143
rect 724 141 726 143
rect 720 140 726 141
rect 731 143 735 145
rect 731 141 732 143
rect 734 141 735 143
rect 731 136 735 141
rect 740 141 746 150
rect 786 149 788 151
rect 790 149 792 151
rect 786 148 792 149
rect 740 139 742 141
rect 744 139 746 141
rect 740 138 746 139
rect 794 144 811 145
rect 794 142 807 144
rect 809 142 811 144
rect 794 141 811 142
rect 825 142 831 151
rect 731 134 732 136
rect 734 135 735 136
rect 734 134 748 135
rect 731 131 748 134
rect 684 129 707 130
rect 684 127 703 129
rect 705 127 707 129
rect 684 126 707 127
rect 664 122 668 124
rect 663 120 668 122
rect 684 120 688 126
rect 663 118 664 120
rect 666 118 668 120
rect 663 116 668 118
rect 672 119 688 120
rect 672 117 674 119
rect 676 117 688 119
rect 672 116 688 117
rect 664 112 668 116
rect 703 120 707 126
rect 703 116 714 120
rect 664 108 688 112
rect 684 105 688 108
rect 710 110 714 116
rect 710 108 711 110
rect 713 108 714 110
rect 710 106 714 108
rect 744 119 748 131
rect 744 117 745 119
rect 747 117 748 119
rect 744 112 748 117
rect 736 108 748 112
rect 684 103 685 105
rect 687 103 688 105
rect 736 104 740 108
rect 751 105 752 107
rect 779 130 780 141
rect 794 137 798 141
rect 825 140 827 142
rect 829 140 831 142
rect 825 139 831 140
rect 836 144 840 146
rect 836 142 837 144
rect 839 142 840 144
rect 783 133 798 137
rect 783 120 787 133
rect 836 137 840 142
rect 845 144 851 151
rect 875 149 876 151
rect 878 149 879 151
rect 845 142 847 144
rect 849 142 851 144
rect 845 141 851 142
rect 875 144 879 149
rect 875 142 876 144
rect 878 142 879 144
rect 875 140 879 142
rect 883 145 916 146
rect 883 143 912 145
rect 914 143 916 145
rect 883 142 916 143
rect 930 142 936 151
rect 836 136 837 137
rect 823 135 837 136
rect 839 135 840 137
rect 823 132 840 135
rect 802 124 808 125
rect 783 118 784 120
rect 786 118 787 120
rect 783 112 787 118
rect 783 111 801 112
rect 783 109 797 111
rect 799 109 801 111
rect 783 108 801 109
rect 720 103 740 104
rect 684 101 688 103
rect 695 102 701 103
rect 695 100 697 102
rect 699 100 701 102
rect 720 101 722 103
rect 724 101 740 103
rect 720 100 740 101
rect 695 94 701 100
rect 823 120 827 132
rect 883 131 887 142
rect 930 140 932 142
rect 934 140 936 142
rect 930 139 936 140
rect 941 144 945 146
rect 941 142 942 144
rect 944 142 945 144
rect 864 130 887 131
rect 864 128 866 130
rect 868 128 887 130
rect 864 127 887 128
rect 864 121 868 127
rect 823 118 824 120
rect 826 118 827 120
rect 823 113 827 118
rect 823 109 835 113
rect 819 106 820 108
rect 831 105 835 109
rect 857 117 868 121
rect 857 111 861 117
rect 883 121 887 127
rect 891 137 895 139
rect 891 135 892 137
rect 894 135 895 137
rect 891 130 895 135
rect 891 128 892 130
rect 894 129 895 130
rect 894 128 907 129
rect 891 125 907 128
rect 903 123 907 125
rect 903 121 908 123
rect 883 120 899 121
rect 883 118 895 120
rect 897 118 899 120
rect 883 117 899 118
rect 903 119 905 121
rect 907 119 908 121
rect 903 117 908 119
rect 857 109 858 111
rect 860 109 861 111
rect 857 107 861 109
rect 903 113 907 117
rect 883 109 907 113
rect 883 106 887 109
rect 831 104 851 105
rect 883 104 884 106
rect 886 104 887 106
rect 831 102 847 104
rect 849 102 851 104
rect 831 101 851 102
rect 870 103 876 104
rect 870 101 872 103
rect 874 101 876 103
rect 883 102 887 104
rect 941 137 945 142
rect 950 144 956 151
rect 980 149 981 151
rect 983 149 984 151
rect 950 142 952 144
rect 954 142 956 144
rect 950 141 956 142
rect 980 144 984 149
rect 1036 149 1038 151
rect 1040 149 1042 151
rect 1036 148 1042 149
rect 980 142 981 144
rect 983 142 984 144
rect 980 140 984 142
rect 988 145 1021 146
rect 988 143 1017 145
rect 1019 143 1021 145
rect 988 142 1021 143
rect 941 136 942 137
rect 928 135 942 136
rect 944 135 945 137
rect 928 132 945 135
rect 928 120 932 132
rect 988 131 992 142
rect 1044 144 1061 145
rect 1044 142 1057 144
rect 1059 142 1061 144
rect 1044 141 1061 142
rect 1075 142 1081 151
rect 969 130 992 131
rect 969 128 971 130
rect 973 128 992 130
rect 969 127 992 128
rect 969 121 973 127
rect 928 118 929 120
rect 931 118 932 120
rect 928 113 932 118
rect 928 109 940 113
rect 924 106 925 108
rect 786 98 792 99
rect 786 96 788 98
rect 790 96 792 98
rect 786 95 792 96
rect 805 98 811 99
rect 805 96 807 98
rect 809 96 811 98
rect 805 95 811 96
rect 870 95 876 101
rect 936 105 940 109
rect 962 117 973 121
rect 962 111 966 117
rect 988 121 992 127
rect 996 137 1000 139
rect 996 135 997 137
rect 999 135 1000 137
rect 996 130 1000 135
rect 996 128 997 130
rect 999 129 1000 130
rect 999 128 1012 129
rect 996 125 1012 128
rect 1008 123 1012 125
rect 1008 121 1013 123
rect 988 120 1004 121
rect 988 118 1000 120
rect 1002 118 1004 120
rect 988 117 1004 118
rect 1008 119 1010 121
rect 1012 119 1013 121
rect 1008 117 1013 119
rect 962 109 963 111
rect 965 109 966 111
rect 962 107 966 109
rect 1008 113 1012 117
rect 988 109 1012 113
rect 988 106 992 109
rect 936 104 956 105
rect 988 104 989 106
rect 991 104 992 106
rect 1029 130 1030 141
rect 1044 137 1048 141
rect 1075 140 1077 142
rect 1079 140 1081 142
rect 1075 139 1081 140
rect 1086 144 1090 146
rect 1086 142 1087 144
rect 1089 142 1090 144
rect 1033 133 1048 137
rect 1033 120 1037 133
rect 1086 137 1090 142
rect 1095 144 1101 151
rect 1125 149 1126 151
rect 1128 149 1129 151
rect 1095 142 1097 144
rect 1099 142 1101 144
rect 1095 141 1101 142
rect 1125 144 1129 149
rect 1125 142 1126 144
rect 1128 142 1129 144
rect 1125 140 1129 142
rect 1133 145 1166 146
rect 1133 143 1162 145
rect 1164 143 1166 145
rect 1133 142 1166 143
rect 1180 142 1186 151
rect 1086 136 1087 137
rect 1073 135 1087 136
rect 1089 135 1090 137
rect 1073 132 1090 135
rect 1052 124 1058 125
rect 1033 118 1034 120
rect 1036 118 1037 120
rect 1033 112 1037 118
rect 1033 111 1051 112
rect 1033 109 1047 111
rect 1049 109 1051 111
rect 1033 108 1051 109
rect 936 102 952 104
rect 954 102 956 104
rect 936 101 956 102
rect 975 103 981 104
rect 975 101 977 103
rect 979 101 981 103
rect 988 102 992 104
rect 1073 120 1077 132
rect 1133 131 1137 142
rect 1180 140 1182 142
rect 1184 140 1186 142
rect 1180 139 1186 140
rect 1191 144 1195 146
rect 1191 142 1192 144
rect 1194 142 1195 144
rect 1114 130 1137 131
rect 1114 128 1116 130
rect 1118 128 1137 130
rect 1114 127 1137 128
rect 1114 121 1118 127
rect 1073 118 1074 120
rect 1076 118 1077 120
rect 1073 113 1077 118
rect 1073 109 1085 113
rect 1069 106 1070 108
rect 975 95 981 101
rect 1081 105 1085 109
rect 1107 117 1118 121
rect 1107 111 1111 117
rect 1133 121 1137 127
rect 1141 137 1145 139
rect 1141 135 1142 137
rect 1144 135 1145 137
rect 1141 130 1145 135
rect 1141 128 1142 130
rect 1144 129 1145 130
rect 1144 128 1157 129
rect 1141 125 1157 128
rect 1153 123 1157 125
rect 1153 121 1158 123
rect 1133 120 1149 121
rect 1133 118 1145 120
rect 1147 118 1149 120
rect 1133 117 1149 118
rect 1153 119 1155 121
rect 1157 119 1158 121
rect 1153 117 1158 119
rect 1107 109 1108 111
rect 1110 109 1111 111
rect 1107 107 1111 109
rect 1153 113 1157 117
rect 1133 109 1157 113
rect 1133 106 1137 109
rect 1081 104 1101 105
rect 1133 104 1134 106
rect 1136 104 1137 106
rect 1081 102 1097 104
rect 1099 102 1101 104
rect 1081 101 1101 102
rect 1120 103 1126 104
rect 1120 101 1122 103
rect 1124 101 1126 103
rect 1133 102 1137 104
rect 1191 137 1195 142
rect 1200 144 1206 151
rect 1230 149 1231 151
rect 1233 149 1234 151
rect 1200 142 1202 144
rect 1204 142 1206 144
rect 1200 141 1206 142
rect 1230 144 1234 149
rect 1286 149 1288 151
rect 1290 149 1292 151
rect 1286 148 1292 149
rect 1230 142 1231 144
rect 1233 142 1234 144
rect 1230 140 1234 142
rect 1238 145 1271 146
rect 1238 143 1267 145
rect 1269 143 1271 145
rect 1238 142 1271 143
rect 1191 136 1192 137
rect 1178 135 1192 136
rect 1194 135 1195 137
rect 1178 132 1195 135
rect 1178 120 1182 132
rect 1238 131 1242 142
rect 1294 144 1311 145
rect 1294 142 1307 144
rect 1309 142 1311 144
rect 1294 141 1311 142
rect 1325 142 1331 151
rect 1219 130 1242 131
rect 1219 128 1221 130
rect 1223 128 1242 130
rect 1219 127 1242 128
rect 1219 121 1223 127
rect 1178 118 1179 120
rect 1181 118 1182 120
rect 1178 113 1182 118
rect 1178 109 1190 113
rect 1174 106 1175 108
rect 1036 98 1042 99
rect 1036 96 1038 98
rect 1040 96 1042 98
rect 1036 95 1042 96
rect 1055 98 1061 99
rect 1055 96 1057 98
rect 1059 96 1061 98
rect 1055 95 1061 96
rect 1120 95 1126 101
rect 1186 105 1190 109
rect 1212 117 1223 121
rect 1212 111 1216 117
rect 1238 121 1242 127
rect 1246 137 1250 139
rect 1246 135 1247 137
rect 1249 135 1250 137
rect 1246 130 1250 135
rect 1246 128 1247 130
rect 1249 129 1250 130
rect 1249 128 1262 129
rect 1246 125 1262 128
rect 1258 123 1262 125
rect 1258 121 1263 123
rect 1238 120 1254 121
rect 1238 118 1250 120
rect 1252 118 1254 120
rect 1238 117 1254 118
rect 1258 119 1260 121
rect 1262 119 1263 121
rect 1258 117 1263 119
rect 1212 109 1213 111
rect 1215 109 1216 111
rect 1212 107 1216 109
rect 1258 113 1262 117
rect 1238 109 1262 113
rect 1238 106 1242 109
rect 1186 104 1206 105
rect 1238 104 1239 106
rect 1241 104 1242 106
rect 1279 130 1280 141
rect 1294 137 1298 141
rect 1325 140 1327 142
rect 1329 140 1331 142
rect 1325 139 1331 140
rect 1336 144 1340 146
rect 1336 142 1337 144
rect 1339 142 1340 144
rect 1283 133 1298 137
rect 1283 120 1287 133
rect 1336 137 1340 142
rect 1345 144 1351 151
rect 1375 149 1376 151
rect 1378 149 1379 151
rect 1345 142 1347 144
rect 1349 142 1351 144
rect 1345 141 1351 142
rect 1375 144 1379 149
rect 1375 142 1376 144
rect 1378 142 1379 144
rect 1375 140 1379 142
rect 1383 145 1416 146
rect 1383 143 1412 145
rect 1414 143 1416 145
rect 1383 142 1416 143
rect 1430 142 1436 151
rect 1336 136 1337 137
rect 1323 135 1337 136
rect 1339 135 1340 137
rect 1323 132 1340 135
rect 1302 124 1308 125
rect 1283 118 1284 120
rect 1286 118 1287 120
rect 1283 112 1287 118
rect 1283 111 1301 112
rect 1283 109 1297 111
rect 1299 109 1301 111
rect 1283 108 1301 109
rect 1186 102 1202 104
rect 1204 102 1206 104
rect 1186 101 1206 102
rect 1225 103 1231 104
rect 1225 101 1227 103
rect 1229 101 1231 103
rect 1238 102 1242 104
rect 1323 120 1327 132
rect 1383 131 1387 142
rect 1430 140 1432 142
rect 1434 140 1436 142
rect 1430 139 1436 140
rect 1441 144 1445 146
rect 1441 142 1442 144
rect 1444 142 1445 144
rect 1364 130 1387 131
rect 1364 128 1366 130
rect 1368 128 1387 130
rect 1364 127 1387 128
rect 1364 121 1368 127
rect 1323 118 1324 120
rect 1326 118 1327 120
rect 1323 113 1327 118
rect 1323 109 1335 113
rect 1319 106 1320 108
rect 1225 95 1231 101
rect 1331 105 1335 109
rect 1357 117 1368 121
rect 1357 111 1361 117
rect 1383 121 1387 127
rect 1391 137 1395 139
rect 1391 135 1392 137
rect 1394 135 1395 137
rect 1391 130 1395 135
rect 1391 128 1392 130
rect 1394 129 1395 130
rect 1394 128 1407 129
rect 1391 125 1407 128
rect 1403 123 1407 125
rect 1403 121 1408 123
rect 1383 120 1399 121
rect 1383 118 1395 120
rect 1397 118 1399 120
rect 1383 117 1399 118
rect 1403 119 1405 121
rect 1407 119 1408 121
rect 1403 117 1408 119
rect 1357 109 1358 111
rect 1360 109 1361 111
rect 1357 107 1361 109
rect 1403 113 1407 117
rect 1383 109 1407 113
rect 1383 106 1387 109
rect 1331 104 1351 105
rect 1383 104 1384 106
rect 1386 104 1387 106
rect 1331 102 1347 104
rect 1349 102 1351 104
rect 1331 101 1351 102
rect 1370 103 1376 104
rect 1370 101 1372 103
rect 1374 101 1376 103
rect 1383 102 1387 104
rect 1441 137 1445 142
rect 1450 144 1456 151
rect 1480 149 1481 151
rect 1483 149 1484 151
rect 1450 142 1452 144
rect 1454 142 1456 144
rect 1450 141 1456 142
rect 1480 144 1484 149
rect 1536 149 1538 151
rect 1540 149 1542 151
rect 1536 148 1542 149
rect 1480 142 1481 144
rect 1483 142 1484 144
rect 1480 140 1484 142
rect 1488 145 1521 146
rect 1488 143 1517 145
rect 1519 143 1521 145
rect 1488 142 1521 143
rect 1441 136 1442 137
rect 1428 135 1442 136
rect 1444 135 1445 137
rect 1428 132 1445 135
rect 1428 120 1432 132
rect 1488 131 1492 142
rect 1544 144 1561 145
rect 1544 142 1557 144
rect 1559 142 1561 144
rect 1544 141 1561 142
rect 1575 142 1581 151
rect 1469 130 1492 131
rect 1469 128 1471 130
rect 1473 128 1492 130
rect 1469 127 1492 128
rect 1469 121 1473 127
rect 1428 118 1429 120
rect 1431 118 1432 120
rect 1428 113 1432 118
rect 1428 109 1440 113
rect 1424 106 1425 108
rect 1286 98 1292 99
rect 1286 96 1288 98
rect 1290 96 1292 98
rect 1286 95 1292 96
rect 1305 98 1311 99
rect 1305 96 1307 98
rect 1309 96 1311 98
rect 1305 95 1311 96
rect 1370 95 1376 101
rect 1436 105 1440 109
rect 1462 117 1473 121
rect 1462 111 1466 117
rect 1488 121 1492 127
rect 1496 137 1500 139
rect 1496 135 1497 137
rect 1499 135 1500 137
rect 1496 130 1500 135
rect 1496 128 1497 130
rect 1499 129 1500 130
rect 1499 128 1512 129
rect 1496 125 1512 128
rect 1508 123 1512 125
rect 1508 121 1513 123
rect 1488 120 1504 121
rect 1488 118 1500 120
rect 1502 118 1504 120
rect 1488 117 1504 118
rect 1508 119 1510 121
rect 1512 119 1513 121
rect 1508 117 1513 119
rect 1462 109 1463 111
rect 1465 109 1466 111
rect 1462 107 1466 109
rect 1508 113 1512 117
rect 1488 109 1512 113
rect 1488 106 1492 109
rect 1436 104 1456 105
rect 1488 104 1489 106
rect 1491 104 1492 106
rect 1529 130 1530 141
rect 1544 137 1548 141
rect 1575 140 1577 142
rect 1579 140 1581 142
rect 1575 139 1581 140
rect 1586 144 1590 146
rect 1586 142 1587 144
rect 1589 142 1590 144
rect 1533 133 1548 137
rect 1533 120 1537 133
rect 1586 137 1590 142
rect 1595 144 1601 151
rect 1625 149 1626 151
rect 1628 149 1629 151
rect 1595 142 1597 144
rect 1599 142 1601 144
rect 1595 141 1601 142
rect 1625 144 1629 149
rect 1625 142 1626 144
rect 1628 142 1629 144
rect 1625 140 1629 142
rect 1633 145 1666 146
rect 1633 143 1662 145
rect 1664 143 1666 145
rect 1633 142 1666 143
rect 1680 142 1686 151
rect 1586 136 1587 137
rect 1573 135 1587 136
rect 1589 135 1590 137
rect 1573 132 1590 135
rect 1552 124 1558 125
rect 1533 118 1534 120
rect 1536 118 1537 120
rect 1533 112 1537 118
rect 1533 111 1551 112
rect 1533 109 1547 111
rect 1549 109 1551 111
rect 1533 108 1551 109
rect 1436 102 1452 104
rect 1454 102 1456 104
rect 1436 101 1456 102
rect 1475 103 1481 104
rect 1475 101 1477 103
rect 1479 101 1481 103
rect 1488 102 1492 104
rect 1573 120 1577 132
rect 1633 131 1637 142
rect 1680 140 1682 142
rect 1684 140 1686 142
rect 1680 139 1686 140
rect 1691 144 1695 146
rect 1691 142 1692 144
rect 1694 142 1695 144
rect 1614 130 1637 131
rect 1614 128 1616 130
rect 1618 128 1637 130
rect 1614 127 1637 128
rect 1614 121 1618 127
rect 1573 118 1574 120
rect 1576 118 1577 120
rect 1573 113 1577 118
rect 1573 109 1585 113
rect 1569 106 1570 108
rect 1475 95 1481 101
rect 1581 105 1585 109
rect 1607 117 1618 121
rect 1607 111 1611 117
rect 1633 121 1637 127
rect 1641 137 1645 139
rect 1641 135 1642 137
rect 1644 135 1645 137
rect 1641 130 1645 135
rect 1641 128 1642 130
rect 1644 129 1645 130
rect 1644 128 1657 129
rect 1641 125 1657 128
rect 1653 123 1657 125
rect 1653 121 1658 123
rect 1633 120 1649 121
rect 1633 118 1645 120
rect 1647 118 1649 120
rect 1633 117 1649 118
rect 1653 119 1655 121
rect 1657 119 1658 121
rect 1653 117 1658 119
rect 1607 109 1608 111
rect 1610 109 1611 111
rect 1607 107 1611 109
rect 1653 113 1657 117
rect 1633 109 1657 113
rect 1633 106 1637 109
rect 1581 104 1601 105
rect 1633 104 1634 106
rect 1636 104 1637 106
rect 1581 102 1597 104
rect 1599 102 1601 104
rect 1581 101 1601 102
rect 1620 103 1626 104
rect 1620 101 1622 103
rect 1624 101 1626 103
rect 1633 102 1637 104
rect 1691 137 1695 142
rect 1700 144 1706 151
rect 1730 149 1731 151
rect 1733 149 1734 151
rect 1700 142 1702 144
rect 1704 142 1706 144
rect 1700 141 1706 142
rect 1730 144 1734 149
rect 1730 142 1731 144
rect 1733 142 1734 144
rect 1730 140 1734 142
rect 1738 145 1771 146
rect 1738 143 1767 145
rect 1769 143 1771 145
rect 1738 142 1771 143
rect 1833 142 1839 151
rect 1691 136 1692 137
rect 1678 135 1692 136
rect 1694 135 1695 137
rect 1678 132 1695 135
rect 1678 120 1682 132
rect 1738 131 1742 142
rect 1833 140 1835 142
rect 1837 140 1839 142
rect 1833 139 1839 140
rect 1844 144 1848 146
rect 1844 142 1845 144
rect 1847 142 1848 144
rect 1719 130 1742 131
rect 1719 128 1721 130
rect 1723 128 1742 130
rect 1719 127 1742 128
rect 1719 121 1723 127
rect 1678 118 1679 120
rect 1681 118 1682 120
rect 1678 113 1682 118
rect 1678 109 1690 113
rect 1674 106 1675 108
rect 1536 98 1542 99
rect 1536 96 1538 98
rect 1540 96 1542 98
rect 1536 95 1542 96
rect 1555 98 1561 99
rect 1555 96 1557 98
rect 1559 96 1561 98
rect 1555 95 1561 96
rect 1620 95 1626 101
rect 1686 105 1690 109
rect 1712 117 1723 121
rect 1712 111 1716 117
rect 1738 121 1742 127
rect 1746 137 1750 139
rect 1746 135 1747 137
rect 1749 135 1750 137
rect 1746 130 1750 135
rect 1746 128 1747 130
rect 1749 129 1750 130
rect 1749 128 1762 129
rect 1746 125 1762 128
rect 1758 123 1762 125
rect 1758 121 1763 123
rect 1738 120 1754 121
rect 1738 118 1750 120
rect 1752 118 1754 120
rect 1738 117 1754 118
rect 1758 119 1760 121
rect 1762 119 1763 121
rect 1758 117 1763 119
rect 1712 109 1713 111
rect 1715 109 1716 111
rect 1712 107 1716 109
rect 1758 113 1762 117
rect 1738 109 1762 113
rect 1738 106 1742 109
rect 1686 104 1706 105
rect 1738 104 1739 106
rect 1741 104 1742 106
rect 1686 102 1702 104
rect 1704 102 1706 104
rect 1686 101 1706 102
rect 1725 103 1731 104
rect 1725 101 1727 103
rect 1729 101 1731 103
rect 1738 102 1742 104
rect 1844 137 1848 142
rect 1853 144 1859 151
rect 1853 142 1855 144
rect 1857 142 1859 144
rect 1853 141 1859 142
rect 1863 144 1869 151
rect 1863 142 1865 144
rect 1867 142 1869 144
rect 1863 141 1869 142
rect 1874 144 1878 146
rect 1874 142 1875 144
rect 1877 142 1878 144
rect 1844 136 1845 137
rect 1831 135 1845 136
rect 1847 135 1848 137
rect 1831 132 1848 135
rect 1831 120 1835 132
rect 1874 137 1878 142
rect 1883 142 1889 151
rect 1883 140 1885 142
rect 1887 140 1889 142
rect 1883 139 1889 140
rect 1913 142 1919 151
rect 1913 140 1915 142
rect 1917 140 1919 142
rect 1913 139 1919 140
rect 1924 144 1928 146
rect 1924 142 1925 144
rect 1927 142 1928 144
rect 1874 135 1875 137
rect 1877 136 1878 137
rect 1877 135 1891 136
rect 1874 132 1891 135
rect 1831 118 1832 120
rect 1834 118 1835 120
rect 1831 113 1835 118
rect 1831 109 1843 113
rect 1827 106 1828 108
rect 1725 95 1731 101
rect 1839 105 1843 109
rect 1887 120 1891 132
rect 1887 118 1888 120
rect 1890 118 1891 120
rect 1887 113 1891 118
rect 1879 109 1891 113
rect 1879 105 1883 109
rect 1894 106 1895 108
rect 1839 104 1859 105
rect 1839 102 1855 104
rect 1857 102 1859 104
rect 1839 101 1859 102
rect 1863 104 1883 105
rect 1863 102 1865 104
rect 1867 102 1883 104
rect 1863 101 1883 102
rect 1924 137 1928 142
rect 1933 144 1939 151
rect 1963 149 1964 151
rect 1966 149 1967 151
rect 1933 142 1935 144
rect 1937 142 1939 144
rect 1933 141 1939 142
rect 1963 144 1967 149
rect 1963 142 1964 144
rect 1966 142 1967 144
rect 1963 140 1967 142
rect 1971 145 2004 146
rect 1971 143 2000 145
rect 2002 143 2004 145
rect 1971 142 2004 143
rect 1924 136 1925 137
rect 1911 135 1925 136
rect 1927 135 1928 137
rect 1911 132 1928 135
rect 1911 120 1915 132
rect 1971 131 1975 142
rect 1952 130 1975 131
rect 1952 128 1954 130
rect 1956 128 1975 130
rect 1952 127 1975 128
rect 1952 121 1956 127
rect 1911 118 1912 120
rect 1914 118 1915 120
rect 1911 113 1915 118
rect 1911 109 1923 113
rect 1907 106 1908 108
rect 1919 105 1923 109
rect 1945 117 1956 121
rect 1945 111 1949 117
rect 1971 121 1975 127
rect 1979 137 1983 139
rect 1979 135 1980 137
rect 1982 135 1983 137
rect 1979 130 1983 135
rect 1979 128 1980 130
rect 1982 129 1983 130
rect 1982 128 1995 129
rect 1979 125 1995 128
rect 1991 123 1995 125
rect 1991 121 1996 123
rect 1971 120 1987 121
rect 1971 118 1983 120
rect 1985 118 1987 120
rect 1971 117 1987 118
rect 1991 119 1993 121
rect 1995 119 1996 121
rect 1991 117 1996 119
rect 1945 109 1946 111
rect 1948 109 1949 111
rect 1945 107 1949 109
rect 1991 113 1995 117
rect 1971 109 1995 113
rect 1971 106 1975 109
rect 1919 104 1939 105
rect 1971 104 1972 106
rect 1974 104 1975 106
rect 1919 102 1935 104
rect 1937 102 1939 104
rect 1919 101 1939 102
rect 1958 103 1964 104
rect 1958 101 1960 103
rect 1962 101 1964 103
rect 1971 102 1975 104
rect 1958 95 1964 101
rect 18 68 24 69
rect 18 66 20 68
rect 22 66 24 68
rect 18 65 24 66
rect 37 68 43 69
rect 37 66 39 68
rect 41 66 43 68
rect 37 65 43 66
rect 102 63 108 69
rect 63 62 83 63
rect 63 60 79 62
rect 81 60 83 62
rect 102 61 104 63
rect 106 61 108 63
rect 102 60 108 61
rect 115 60 119 62
rect 63 59 83 60
rect 15 55 33 56
rect 15 53 29 55
rect 31 53 33 55
rect 15 52 33 53
rect 15 46 19 52
rect 51 56 52 58
rect 63 55 67 59
rect 115 58 116 60
rect 118 58 119 60
rect 15 44 16 46
rect 18 44 19 46
rect 11 23 12 34
rect 15 31 19 44
rect 34 39 40 40
rect 15 27 30 31
rect 26 23 30 27
rect 55 51 67 55
rect 55 46 59 51
rect 55 44 56 46
rect 58 44 59 46
rect 55 32 59 44
rect 89 55 93 57
rect 89 53 90 55
rect 92 53 93 55
rect 89 47 93 53
rect 115 55 119 58
rect 115 51 139 55
rect 89 43 100 47
rect 96 37 100 43
rect 135 47 139 51
rect 115 46 131 47
rect 115 44 127 46
rect 129 44 131 46
rect 115 43 131 44
rect 135 45 140 47
rect 135 43 137 45
rect 139 43 140 45
rect 115 37 119 43
rect 135 41 140 43
rect 135 39 139 41
rect 96 36 119 37
rect 96 34 98 36
rect 100 34 119 36
rect 96 33 119 34
rect 55 29 72 32
rect 55 28 69 29
rect 68 27 69 28
rect 71 27 72 29
rect 57 24 63 25
rect 26 22 43 23
rect 26 20 39 22
rect 41 20 43 22
rect 26 19 43 20
rect 57 22 59 24
rect 61 22 63 24
rect 18 15 24 16
rect 18 13 20 15
rect 22 13 24 15
rect 57 13 63 22
rect 68 22 72 27
rect 68 20 69 22
rect 71 20 72 22
rect 68 18 72 20
rect 77 22 83 23
rect 77 20 79 22
rect 81 20 83 22
rect 77 13 83 20
rect 107 22 111 24
rect 107 20 108 22
rect 110 20 111 22
rect 107 15 111 20
rect 115 22 119 33
rect 123 36 139 39
rect 123 34 124 36
rect 126 35 139 36
rect 126 34 127 35
rect 123 29 127 34
rect 123 27 124 29
rect 126 27 127 29
rect 123 25 127 27
rect 207 63 213 69
rect 268 68 274 69
rect 268 66 270 68
rect 272 66 274 68
rect 268 65 274 66
rect 287 68 293 69
rect 287 66 289 68
rect 291 66 293 68
rect 287 65 293 66
rect 168 62 188 63
rect 168 60 184 62
rect 186 60 188 62
rect 207 61 209 63
rect 211 61 213 63
rect 207 60 213 61
rect 220 60 224 62
rect 168 59 188 60
rect 156 56 157 58
rect 168 55 172 59
rect 220 58 221 60
rect 223 58 224 60
rect 160 51 172 55
rect 160 46 164 51
rect 160 44 161 46
rect 163 44 164 46
rect 160 32 164 44
rect 194 55 198 57
rect 194 53 195 55
rect 197 53 198 55
rect 194 47 198 53
rect 220 55 224 58
rect 220 51 244 55
rect 194 43 205 47
rect 201 37 205 43
rect 240 47 244 51
rect 220 46 236 47
rect 220 44 232 46
rect 234 44 236 46
rect 220 43 236 44
rect 240 45 245 47
rect 240 43 242 45
rect 244 43 245 45
rect 220 37 224 43
rect 240 41 245 43
rect 240 39 244 41
rect 201 36 224 37
rect 201 34 203 36
rect 205 34 224 36
rect 201 33 224 34
rect 160 29 177 32
rect 160 28 174 29
rect 173 27 174 28
rect 176 27 177 29
rect 162 24 168 25
rect 162 22 164 24
rect 166 22 168 24
rect 115 21 148 22
rect 115 19 144 21
rect 146 19 148 21
rect 115 18 148 19
rect 107 13 108 15
rect 110 13 111 15
rect 162 13 168 22
rect 173 22 177 27
rect 173 20 174 22
rect 176 20 177 22
rect 173 18 177 20
rect 182 22 188 23
rect 182 20 184 22
rect 186 20 188 22
rect 182 13 188 20
rect 212 22 216 24
rect 212 20 213 22
rect 215 20 216 22
rect 212 15 216 20
rect 220 22 224 33
rect 228 36 244 39
rect 228 34 229 36
rect 231 35 244 36
rect 231 34 232 35
rect 228 29 232 34
rect 352 63 358 69
rect 313 62 333 63
rect 313 60 329 62
rect 331 60 333 62
rect 352 61 354 63
rect 356 61 358 63
rect 352 60 358 61
rect 365 60 369 62
rect 313 59 333 60
rect 228 27 229 29
rect 231 27 232 29
rect 228 25 232 27
rect 265 55 283 56
rect 265 53 279 55
rect 281 53 283 55
rect 265 52 283 53
rect 265 46 269 52
rect 301 56 302 58
rect 313 55 317 59
rect 365 58 366 60
rect 368 58 369 60
rect 265 44 266 46
rect 268 44 269 46
rect 261 23 262 34
rect 265 31 269 44
rect 284 39 290 40
rect 265 27 280 31
rect 276 23 280 27
rect 305 51 317 55
rect 305 46 309 51
rect 305 44 306 46
rect 308 44 309 46
rect 305 32 309 44
rect 339 55 343 57
rect 339 53 340 55
rect 342 53 343 55
rect 339 47 343 53
rect 365 55 369 58
rect 365 51 389 55
rect 339 43 350 47
rect 346 37 350 43
rect 385 47 389 51
rect 365 46 381 47
rect 365 44 377 46
rect 379 44 381 46
rect 365 43 381 44
rect 385 45 390 47
rect 385 43 387 45
rect 389 43 390 45
rect 365 37 369 43
rect 385 41 390 43
rect 385 39 389 41
rect 346 36 369 37
rect 346 34 348 36
rect 350 34 369 36
rect 346 33 369 34
rect 305 29 322 32
rect 305 28 319 29
rect 318 27 319 28
rect 321 27 322 29
rect 307 24 313 25
rect 220 21 253 22
rect 220 19 249 21
rect 251 19 253 21
rect 220 18 253 19
rect 276 22 293 23
rect 276 20 289 22
rect 291 20 293 22
rect 276 19 293 20
rect 307 22 309 24
rect 311 22 313 24
rect 212 13 213 15
rect 215 13 216 15
rect 268 15 274 16
rect 268 13 270 15
rect 272 13 274 15
rect 307 13 313 22
rect 318 22 322 27
rect 318 20 319 22
rect 321 20 322 22
rect 318 18 322 20
rect 327 22 333 23
rect 327 20 329 22
rect 331 20 333 22
rect 327 13 333 20
rect 357 22 361 24
rect 357 20 358 22
rect 360 20 361 22
rect 357 15 361 20
rect 365 22 369 33
rect 373 36 389 39
rect 373 34 374 36
rect 376 35 389 36
rect 376 34 377 35
rect 373 29 377 34
rect 373 27 374 29
rect 376 27 377 29
rect 373 25 377 27
rect 457 63 463 69
rect 518 68 524 69
rect 518 66 520 68
rect 522 66 524 68
rect 518 65 524 66
rect 537 68 543 69
rect 537 66 539 68
rect 541 66 543 68
rect 537 65 543 66
rect 418 62 438 63
rect 418 60 434 62
rect 436 60 438 62
rect 457 61 459 63
rect 461 61 463 63
rect 457 60 463 61
rect 470 60 474 62
rect 418 59 438 60
rect 406 56 407 58
rect 418 55 422 59
rect 470 58 471 60
rect 473 58 474 60
rect 410 51 422 55
rect 410 46 414 51
rect 410 44 411 46
rect 413 44 414 46
rect 410 32 414 44
rect 444 55 448 57
rect 444 53 445 55
rect 447 53 448 55
rect 444 47 448 53
rect 470 55 474 58
rect 470 51 494 55
rect 444 43 455 47
rect 451 37 455 43
rect 490 47 494 51
rect 470 46 486 47
rect 470 44 482 46
rect 484 44 486 46
rect 470 43 486 44
rect 490 45 495 47
rect 490 43 492 45
rect 494 43 495 45
rect 470 37 474 43
rect 490 41 495 43
rect 490 39 494 41
rect 451 36 474 37
rect 451 34 453 36
rect 455 34 474 36
rect 451 33 474 34
rect 410 29 427 32
rect 410 28 424 29
rect 423 27 424 28
rect 426 27 427 29
rect 412 24 418 25
rect 412 22 414 24
rect 416 22 418 24
rect 365 21 398 22
rect 365 19 394 21
rect 396 19 398 21
rect 365 18 398 19
rect 357 13 358 15
rect 360 13 361 15
rect 412 13 418 22
rect 423 22 427 27
rect 423 20 424 22
rect 426 20 427 22
rect 423 18 427 20
rect 432 22 438 23
rect 432 20 434 22
rect 436 20 438 22
rect 432 13 438 20
rect 462 22 466 24
rect 462 20 463 22
rect 465 20 466 22
rect 462 15 466 20
rect 470 22 474 33
rect 478 36 494 39
rect 478 34 479 36
rect 481 35 494 36
rect 481 34 482 35
rect 478 29 482 34
rect 602 63 608 69
rect 563 62 583 63
rect 563 60 579 62
rect 581 60 583 62
rect 602 61 604 63
rect 606 61 608 63
rect 602 60 608 61
rect 615 60 619 62
rect 563 59 583 60
rect 478 27 479 29
rect 481 27 482 29
rect 478 25 482 27
rect 515 55 533 56
rect 515 53 529 55
rect 531 53 533 55
rect 515 52 533 53
rect 515 46 519 52
rect 551 56 552 58
rect 563 55 567 59
rect 615 58 616 60
rect 618 58 619 60
rect 515 44 516 46
rect 518 44 519 46
rect 511 23 512 34
rect 515 31 519 44
rect 534 39 540 40
rect 515 27 530 31
rect 526 23 530 27
rect 555 51 567 55
rect 555 46 559 51
rect 555 44 556 46
rect 558 44 559 46
rect 555 32 559 44
rect 589 55 593 57
rect 589 53 590 55
rect 592 53 593 55
rect 589 47 593 53
rect 615 55 619 58
rect 615 51 639 55
rect 589 43 600 47
rect 596 37 600 43
rect 635 47 639 51
rect 615 46 631 47
rect 615 44 627 46
rect 629 44 631 46
rect 615 43 631 44
rect 635 45 640 47
rect 635 43 637 45
rect 639 43 640 45
rect 615 37 619 43
rect 635 41 640 43
rect 635 39 639 41
rect 596 36 619 37
rect 596 34 598 36
rect 600 34 619 36
rect 596 33 619 34
rect 555 29 572 32
rect 555 28 569 29
rect 568 27 569 28
rect 571 27 572 29
rect 557 24 563 25
rect 470 21 503 22
rect 470 19 499 21
rect 501 19 503 21
rect 470 18 503 19
rect 526 22 543 23
rect 526 20 539 22
rect 541 20 543 22
rect 526 19 543 20
rect 557 22 559 24
rect 561 22 563 24
rect 462 13 463 15
rect 465 13 466 15
rect 518 15 524 16
rect 518 13 520 15
rect 522 13 524 15
rect 557 13 563 22
rect 568 22 572 27
rect 568 20 569 22
rect 571 20 572 22
rect 568 18 572 20
rect 577 22 583 23
rect 577 20 579 22
rect 581 20 583 22
rect 577 13 583 20
rect 607 22 611 24
rect 607 20 608 22
rect 610 20 611 22
rect 607 15 611 20
rect 615 22 619 33
rect 623 36 639 39
rect 623 34 624 36
rect 626 35 639 36
rect 626 34 627 35
rect 623 29 627 34
rect 623 27 624 29
rect 626 27 627 29
rect 623 25 627 27
rect 707 63 713 69
rect 768 68 774 69
rect 768 66 770 68
rect 772 66 774 68
rect 768 65 774 66
rect 787 68 793 69
rect 787 66 789 68
rect 791 66 793 68
rect 787 65 793 66
rect 668 62 688 63
rect 668 60 684 62
rect 686 60 688 62
rect 707 61 709 63
rect 711 61 713 63
rect 707 60 713 61
rect 720 60 724 62
rect 668 59 688 60
rect 656 56 657 58
rect 668 55 672 59
rect 720 58 721 60
rect 723 58 724 60
rect 660 51 672 55
rect 660 46 664 51
rect 660 44 661 46
rect 663 44 664 46
rect 660 32 664 44
rect 694 55 698 57
rect 694 53 695 55
rect 697 53 698 55
rect 694 47 698 53
rect 720 55 724 58
rect 720 51 744 55
rect 694 43 705 47
rect 701 37 705 43
rect 740 47 744 51
rect 720 46 736 47
rect 720 44 732 46
rect 734 44 736 46
rect 720 43 736 44
rect 740 45 745 47
rect 740 43 742 45
rect 744 43 745 45
rect 720 37 724 43
rect 740 41 745 43
rect 740 39 744 41
rect 701 36 724 37
rect 701 34 703 36
rect 705 34 724 36
rect 701 33 724 34
rect 660 29 677 32
rect 660 28 674 29
rect 673 27 674 28
rect 676 27 677 29
rect 662 24 668 25
rect 662 22 664 24
rect 666 22 668 24
rect 615 21 648 22
rect 615 19 644 21
rect 646 19 648 21
rect 615 18 648 19
rect 607 13 608 15
rect 610 13 611 15
rect 662 13 668 22
rect 673 22 677 27
rect 673 20 674 22
rect 676 20 677 22
rect 673 18 677 20
rect 682 22 688 23
rect 682 20 684 22
rect 686 20 688 22
rect 682 13 688 20
rect 712 22 716 24
rect 712 20 713 22
rect 715 20 716 22
rect 712 15 716 20
rect 720 22 724 33
rect 728 36 744 39
rect 728 34 729 36
rect 731 35 744 36
rect 731 34 732 35
rect 728 29 732 34
rect 852 63 858 69
rect 813 62 833 63
rect 813 60 829 62
rect 831 60 833 62
rect 852 61 854 63
rect 856 61 858 63
rect 852 60 858 61
rect 865 60 869 62
rect 813 59 833 60
rect 728 27 729 29
rect 731 27 732 29
rect 728 25 732 27
rect 765 55 783 56
rect 765 53 779 55
rect 781 53 783 55
rect 765 52 783 53
rect 765 46 769 52
rect 801 56 802 58
rect 813 55 817 59
rect 865 58 866 60
rect 868 58 869 60
rect 765 44 766 46
rect 768 44 769 46
rect 761 23 762 34
rect 765 31 769 44
rect 784 39 790 40
rect 765 27 780 31
rect 776 23 780 27
rect 805 51 817 55
rect 805 46 809 51
rect 805 44 806 46
rect 808 44 809 46
rect 805 32 809 44
rect 839 55 843 57
rect 839 53 840 55
rect 842 53 843 55
rect 839 47 843 53
rect 865 55 869 58
rect 865 51 889 55
rect 839 43 850 47
rect 846 37 850 43
rect 885 47 889 51
rect 865 46 881 47
rect 865 44 877 46
rect 879 44 881 46
rect 865 43 881 44
rect 885 45 890 47
rect 885 43 887 45
rect 889 43 890 45
rect 865 37 869 43
rect 885 41 890 43
rect 885 39 889 41
rect 846 36 869 37
rect 846 34 848 36
rect 850 34 869 36
rect 846 33 869 34
rect 805 29 822 32
rect 805 28 819 29
rect 818 27 819 28
rect 821 27 822 29
rect 807 24 813 25
rect 720 21 753 22
rect 720 19 749 21
rect 751 19 753 21
rect 720 18 753 19
rect 776 22 793 23
rect 776 20 789 22
rect 791 20 793 22
rect 776 19 793 20
rect 807 22 809 24
rect 811 22 813 24
rect 712 13 713 15
rect 715 13 716 15
rect 768 15 774 16
rect 768 13 770 15
rect 772 13 774 15
rect 807 13 813 22
rect 818 22 822 27
rect 818 20 819 22
rect 821 20 822 22
rect 818 18 822 20
rect 827 22 833 23
rect 827 20 829 22
rect 831 20 833 22
rect 827 13 833 20
rect 857 22 861 24
rect 857 20 858 22
rect 860 20 861 22
rect 857 15 861 20
rect 865 22 869 33
rect 873 36 889 39
rect 873 34 874 36
rect 876 35 889 36
rect 876 34 877 35
rect 873 29 877 34
rect 873 27 874 29
rect 876 27 877 29
rect 873 25 877 27
rect 957 63 963 69
rect 1028 68 1034 69
rect 1028 66 1030 68
rect 1032 66 1034 68
rect 1028 65 1034 66
rect 1047 68 1053 69
rect 1047 66 1049 68
rect 1051 66 1053 68
rect 1047 65 1053 66
rect 918 62 938 63
rect 918 60 934 62
rect 936 60 938 62
rect 957 61 959 63
rect 961 61 963 63
rect 957 60 963 61
rect 970 60 974 62
rect 918 59 938 60
rect 906 56 907 58
rect 918 55 922 59
rect 970 58 971 60
rect 973 58 974 60
rect 910 51 922 55
rect 910 46 914 51
rect 910 44 911 46
rect 913 44 914 46
rect 910 32 914 44
rect 944 55 948 57
rect 944 53 945 55
rect 947 53 948 55
rect 944 47 948 53
rect 970 55 974 58
rect 970 51 994 55
rect 944 43 955 47
rect 951 37 955 43
rect 990 47 994 51
rect 970 46 986 47
rect 970 44 982 46
rect 984 44 986 46
rect 970 43 986 44
rect 990 45 995 47
rect 990 43 992 45
rect 994 43 995 45
rect 970 37 974 43
rect 990 41 995 43
rect 990 39 994 41
rect 951 36 974 37
rect 951 34 953 36
rect 955 34 974 36
rect 951 33 974 34
rect 910 29 927 32
rect 910 28 924 29
rect 923 27 924 28
rect 926 27 927 29
rect 912 24 918 25
rect 912 22 914 24
rect 916 22 918 24
rect 865 21 898 22
rect 865 19 894 21
rect 896 19 898 21
rect 865 18 898 19
rect 857 13 858 15
rect 860 13 861 15
rect 912 13 918 22
rect 923 22 927 27
rect 923 20 924 22
rect 926 20 927 22
rect 923 18 927 20
rect 932 22 938 23
rect 932 20 934 22
rect 936 20 938 22
rect 932 13 938 20
rect 962 22 966 24
rect 962 20 963 22
rect 965 20 966 22
rect 962 15 966 20
rect 970 22 974 33
rect 978 36 994 39
rect 978 34 979 36
rect 981 35 994 36
rect 981 34 982 35
rect 978 29 982 34
rect 1112 63 1118 69
rect 1073 62 1093 63
rect 1073 60 1089 62
rect 1091 60 1093 62
rect 1112 61 1114 63
rect 1116 61 1118 63
rect 1112 60 1118 61
rect 1125 60 1129 62
rect 1073 59 1093 60
rect 978 27 979 29
rect 981 27 982 29
rect 978 25 982 27
rect 1025 55 1043 56
rect 1025 53 1039 55
rect 1041 53 1043 55
rect 1025 52 1043 53
rect 1025 46 1029 52
rect 1061 56 1062 58
rect 1073 55 1077 59
rect 1125 58 1126 60
rect 1128 58 1129 60
rect 1025 44 1026 46
rect 1028 44 1029 46
rect 1021 23 1022 34
rect 1025 31 1029 44
rect 1044 39 1050 40
rect 1025 27 1040 31
rect 1036 23 1040 27
rect 1065 51 1077 55
rect 1065 46 1069 51
rect 1065 44 1066 46
rect 1068 44 1069 46
rect 1065 32 1069 44
rect 1099 55 1103 57
rect 1099 53 1100 55
rect 1102 53 1103 55
rect 1099 47 1103 53
rect 1125 55 1129 58
rect 1125 51 1149 55
rect 1099 43 1110 47
rect 1106 37 1110 43
rect 1145 47 1149 51
rect 1125 46 1141 47
rect 1125 44 1137 46
rect 1139 44 1141 46
rect 1125 43 1141 44
rect 1145 45 1150 47
rect 1145 43 1147 45
rect 1149 43 1150 45
rect 1125 37 1129 43
rect 1145 41 1150 43
rect 1145 39 1149 41
rect 1106 36 1129 37
rect 1106 34 1108 36
rect 1110 34 1129 36
rect 1106 33 1129 34
rect 1065 29 1082 32
rect 1065 28 1079 29
rect 1078 27 1079 28
rect 1081 27 1082 29
rect 1067 24 1073 25
rect 970 21 1003 22
rect 970 19 999 21
rect 1001 19 1003 21
rect 970 18 1003 19
rect 1036 22 1053 23
rect 1036 20 1049 22
rect 1051 20 1053 22
rect 1036 19 1053 20
rect 1067 22 1069 24
rect 1071 22 1073 24
rect 962 13 963 15
rect 965 13 966 15
rect 1028 15 1034 16
rect 1028 13 1030 15
rect 1032 13 1034 15
rect 1067 13 1073 22
rect 1078 22 1082 27
rect 1078 20 1079 22
rect 1081 20 1082 22
rect 1078 18 1082 20
rect 1087 22 1093 23
rect 1087 20 1089 22
rect 1091 20 1093 22
rect 1087 13 1093 20
rect 1117 22 1121 24
rect 1117 20 1118 22
rect 1120 20 1121 22
rect 1117 15 1121 20
rect 1125 22 1129 33
rect 1133 36 1149 39
rect 1133 34 1134 36
rect 1136 35 1149 36
rect 1136 34 1137 35
rect 1133 29 1137 34
rect 1133 27 1134 29
rect 1136 27 1137 29
rect 1133 25 1137 27
rect 1217 63 1223 69
rect 1278 68 1284 69
rect 1278 66 1280 68
rect 1282 66 1284 68
rect 1278 65 1284 66
rect 1297 68 1303 69
rect 1297 66 1299 68
rect 1301 66 1303 68
rect 1297 65 1303 66
rect 1178 62 1198 63
rect 1178 60 1194 62
rect 1196 60 1198 62
rect 1217 61 1219 63
rect 1221 61 1223 63
rect 1217 60 1223 61
rect 1230 60 1234 62
rect 1178 59 1198 60
rect 1166 56 1167 58
rect 1178 55 1182 59
rect 1230 58 1231 60
rect 1233 58 1234 60
rect 1170 51 1182 55
rect 1170 46 1174 51
rect 1170 44 1171 46
rect 1173 44 1174 46
rect 1170 32 1174 44
rect 1204 55 1208 57
rect 1204 53 1205 55
rect 1207 53 1208 55
rect 1204 47 1208 53
rect 1230 55 1234 58
rect 1230 51 1254 55
rect 1204 43 1215 47
rect 1211 37 1215 43
rect 1250 47 1254 51
rect 1230 46 1246 47
rect 1230 44 1242 46
rect 1244 44 1246 46
rect 1230 43 1246 44
rect 1250 45 1255 47
rect 1250 43 1252 45
rect 1254 43 1255 45
rect 1230 37 1234 43
rect 1250 41 1255 43
rect 1250 39 1254 41
rect 1211 36 1234 37
rect 1211 34 1213 36
rect 1215 34 1234 36
rect 1211 33 1234 34
rect 1170 29 1187 32
rect 1170 28 1184 29
rect 1183 27 1184 28
rect 1186 27 1187 29
rect 1172 24 1178 25
rect 1172 22 1174 24
rect 1176 22 1178 24
rect 1125 21 1158 22
rect 1125 19 1154 21
rect 1156 19 1158 21
rect 1125 18 1158 19
rect 1117 13 1118 15
rect 1120 13 1121 15
rect 1172 13 1178 22
rect 1183 22 1187 27
rect 1183 20 1184 22
rect 1186 20 1187 22
rect 1183 18 1187 20
rect 1192 22 1198 23
rect 1192 20 1194 22
rect 1196 20 1198 22
rect 1192 13 1198 20
rect 1222 22 1226 24
rect 1222 20 1223 22
rect 1225 20 1226 22
rect 1222 15 1226 20
rect 1230 22 1234 33
rect 1238 36 1254 39
rect 1238 34 1239 36
rect 1241 35 1254 36
rect 1241 34 1242 35
rect 1238 29 1242 34
rect 1362 63 1368 69
rect 1323 62 1343 63
rect 1323 60 1339 62
rect 1341 60 1343 62
rect 1362 61 1364 63
rect 1366 61 1368 63
rect 1362 60 1368 61
rect 1375 60 1379 62
rect 1323 59 1343 60
rect 1238 27 1239 29
rect 1241 27 1242 29
rect 1238 25 1242 27
rect 1275 55 1293 56
rect 1275 53 1289 55
rect 1291 53 1293 55
rect 1275 52 1293 53
rect 1275 46 1279 52
rect 1311 56 1312 58
rect 1323 55 1327 59
rect 1375 58 1376 60
rect 1378 58 1379 60
rect 1275 44 1276 46
rect 1278 44 1279 46
rect 1271 23 1272 34
rect 1275 31 1279 44
rect 1294 39 1300 40
rect 1275 27 1290 31
rect 1286 23 1290 27
rect 1315 51 1327 55
rect 1315 46 1319 51
rect 1315 44 1316 46
rect 1318 44 1319 46
rect 1315 32 1319 44
rect 1349 55 1353 57
rect 1349 53 1350 55
rect 1352 53 1353 55
rect 1349 47 1353 53
rect 1375 55 1379 58
rect 1375 51 1399 55
rect 1349 43 1360 47
rect 1356 37 1360 43
rect 1395 47 1399 51
rect 1375 46 1391 47
rect 1375 44 1387 46
rect 1389 44 1391 46
rect 1375 43 1391 44
rect 1395 45 1400 47
rect 1395 43 1397 45
rect 1399 43 1400 45
rect 1375 37 1379 43
rect 1395 41 1400 43
rect 1395 39 1399 41
rect 1356 36 1379 37
rect 1356 34 1358 36
rect 1360 34 1379 36
rect 1356 33 1379 34
rect 1315 29 1332 32
rect 1315 28 1329 29
rect 1328 27 1329 28
rect 1331 27 1332 29
rect 1317 24 1323 25
rect 1230 21 1263 22
rect 1230 19 1259 21
rect 1261 19 1263 21
rect 1230 18 1263 19
rect 1286 22 1303 23
rect 1286 20 1299 22
rect 1301 20 1303 22
rect 1286 19 1303 20
rect 1317 22 1319 24
rect 1321 22 1323 24
rect 1222 13 1223 15
rect 1225 13 1226 15
rect 1278 15 1284 16
rect 1278 13 1280 15
rect 1282 13 1284 15
rect 1317 13 1323 22
rect 1328 22 1332 27
rect 1328 20 1329 22
rect 1331 20 1332 22
rect 1328 18 1332 20
rect 1337 22 1343 23
rect 1337 20 1339 22
rect 1341 20 1343 22
rect 1337 13 1343 20
rect 1367 22 1371 24
rect 1367 20 1368 22
rect 1370 20 1371 22
rect 1367 15 1371 20
rect 1375 22 1379 33
rect 1383 36 1399 39
rect 1383 34 1384 36
rect 1386 35 1399 36
rect 1386 34 1387 35
rect 1383 29 1387 34
rect 1383 27 1384 29
rect 1386 27 1387 29
rect 1383 25 1387 27
rect 1467 63 1473 69
rect 1528 68 1534 69
rect 1528 66 1530 68
rect 1532 66 1534 68
rect 1528 65 1534 66
rect 1547 68 1553 69
rect 1547 66 1549 68
rect 1551 66 1553 68
rect 1547 65 1553 66
rect 1428 62 1448 63
rect 1428 60 1444 62
rect 1446 60 1448 62
rect 1467 61 1469 63
rect 1471 61 1473 63
rect 1467 60 1473 61
rect 1480 60 1484 62
rect 1428 59 1448 60
rect 1416 56 1417 58
rect 1428 55 1432 59
rect 1480 58 1481 60
rect 1483 58 1484 60
rect 1420 51 1432 55
rect 1420 46 1424 51
rect 1420 44 1421 46
rect 1423 44 1424 46
rect 1420 32 1424 44
rect 1454 55 1458 57
rect 1454 53 1455 55
rect 1457 53 1458 55
rect 1454 47 1458 53
rect 1480 55 1484 58
rect 1480 51 1504 55
rect 1454 43 1465 47
rect 1461 37 1465 43
rect 1500 47 1504 51
rect 1480 46 1496 47
rect 1480 44 1492 46
rect 1494 44 1496 46
rect 1480 43 1496 44
rect 1500 45 1505 47
rect 1500 43 1502 45
rect 1504 43 1505 45
rect 1480 37 1484 43
rect 1500 41 1505 43
rect 1612 63 1618 69
rect 1573 62 1593 63
rect 1573 60 1589 62
rect 1591 60 1593 62
rect 1612 61 1614 63
rect 1616 61 1618 63
rect 1612 60 1618 61
rect 1625 60 1629 62
rect 1573 59 1593 60
rect 1500 39 1504 41
rect 1461 36 1484 37
rect 1461 34 1463 36
rect 1465 34 1484 36
rect 1461 33 1484 34
rect 1420 29 1437 32
rect 1420 28 1434 29
rect 1433 27 1434 28
rect 1436 27 1437 29
rect 1422 24 1428 25
rect 1422 22 1424 24
rect 1426 22 1428 24
rect 1375 21 1408 22
rect 1375 19 1404 21
rect 1406 19 1408 21
rect 1375 18 1408 19
rect 1367 13 1368 15
rect 1370 13 1371 15
rect 1422 13 1428 22
rect 1433 22 1437 27
rect 1433 20 1434 22
rect 1436 20 1437 22
rect 1433 18 1437 20
rect 1442 22 1448 23
rect 1442 20 1444 22
rect 1446 20 1448 22
rect 1442 13 1448 20
rect 1472 22 1476 24
rect 1472 20 1473 22
rect 1475 20 1476 22
rect 1472 15 1476 20
rect 1480 22 1484 33
rect 1488 36 1504 39
rect 1488 34 1489 36
rect 1491 35 1504 36
rect 1491 34 1492 35
rect 1488 29 1492 34
rect 1488 27 1489 29
rect 1491 27 1492 29
rect 1488 25 1492 27
rect 1525 55 1543 56
rect 1525 53 1539 55
rect 1541 53 1543 55
rect 1525 52 1543 53
rect 1525 46 1529 52
rect 1561 56 1562 58
rect 1573 55 1577 59
rect 1625 58 1626 60
rect 1628 58 1629 60
rect 1525 44 1526 46
rect 1528 44 1529 46
rect 1521 23 1522 34
rect 1525 31 1529 44
rect 1544 39 1550 40
rect 1525 27 1540 31
rect 1536 23 1540 27
rect 1565 51 1577 55
rect 1565 46 1569 51
rect 1565 44 1566 46
rect 1568 44 1569 46
rect 1565 32 1569 44
rect 1599 55 1603 57
rect 1599 53 1600 55
rect 1602 53 1603 55
rect 1599 47 1603 53
rect 1625 55 1629 58
rect 1625 51 1649 55
rect 1599 43 1610 47
rect 1606 37 1610 43
rect 1645 47 1649 51
rect 1625 46 1641 47
rect 1625 44 1637 46
rect 1639 44 1641 46
rect 1625 43 1641 44
rect 1645 45 1650 47
rect 1645 43 1647 45
rect 1649 43 1650 45
rect 1625 37 1629 43
rect 1645 41 1650 43
rect 1645 39 1649 41
rect 1606 36 1629 37
rect 1606 34 1608 36
rect 1610 34 1629 36
rect 1606 33 1629 34
rect 1565 29 1582 32
rect 1565 28 1579 29
rect 1578 27 1579 28
rect 1581 27 1582 29
rect 1567 24 1573 25
rect 1480 21 1513 22
rect 1480 19 1509 21
rect 1511 19 1513 21
rect 1480 18 1513 19
rect 1536 22 1553 23
rect 1536 20 1549 22
rect 1551 20 1553 22
rect 1536 19 1553 20
rect 1567 22 1569 24
rect 1571 22 1573 24
rect 1472 13 1473 15
rect 1475 13 1476 15
rect 1528 15 1534 16
rect 1528 13 1530 15
rect 1532 13 1534 15
rect 1567 13 1573 22
rect 1578 22 1582 27
rect 1578 20 1579 22
rect 1581 20 1582 22
rect 1578 18 1582 20
rect 1587 22 1593 23
rect 1587 20 1589 22
rect 1591 20 1593 22
rect 1587 13 1593 20
rect 1617 22 1621 24
rect 1617 20 1618 22
rect 1620 20 1621 22
rect 1617 15 1621 20
rect 1625 22 1629 33
rect 1633 36 1649 39
rect 1633 34 1634 36
rect 1636 35 1649 36
rect 1636 34 1637 35
rect 1633 29 1637 34
rect 1633 27 1634 29
rect 1636 27 1637 29
rect 1633 25 1637 27
rect 1717 63 1723 69
rect 1778 68 1784 69
rect 1778 66 1780 68
rect 1782 66 1784 68
rect 1778 65 1784 66
rect 1797 68 1803 69
rect 1797 66 1799 68
rect 1801 66 1803 68
rect 1797 65 1803 66
rect 1678 62 1698 63
rect 1678 60 1694 62
rect 1696 60 1698 62
rect 1717 61 1719 63
rect 1721 61 1723 63
rect 1717 60 1723 61
rect 1730 60 1734 62
rect 1678 59 1698 60
rect 1666 56 1667 58
rect 1678 55 1682 59
rect 1730 58 1731 60
rect 1733 58 1734 60
rect 1670 51 1682 55
rect 1670 46 1674 51
rect 1670 44 1671 46
rect 1673 44 1674 46
rect 1670 32 1674 44
rect 1704 55 1708 57
rect 1704 53 1705 55
rect 1707 53 1708 55
rect 1704 47 1708 53
rect 1730 55 1734 58
rect 1730 51 1754 55
rect 1704 43 1715 47
rect 1711 37 1715 43
rect 1750 47 1754 51
rect 1730 46 1746 47
rect 1730 44 1742 46
rect 1744 44 1746 46
rect 1730 43 1746 44
rect 1750 45 1755 47
rect 1750 43 1752 45
rect 1754 43 1755 45
rect 1730 37 1734 43
rect 1750 41 1755 43
rect 1750 39 1754 41
rect 1711 36 1734 37
rect 1711 34 1713 36
rect 1715 34 1734 36
rect 1711 33 1734 34
rect 1670 29 1687 32
rect 1670 28 1684 29
rect 1683 27 1684 28
rect 1686 27 1687 29
rect 1672 24 1678 25
rect 1672 22 1674 24
rect 1676 22 1678 24
rect 1625 21 1658 22
rect 1625 19 1654 21
rect 1656 19 1658 21
rect 1625 18 1658 19
rect 1617 13 1618 15
rect 1620 13 1621 15
rect 1672 13 1678 22
rect 1683 22 1687 27
rect 1683 20 1684 22
rect 1686 20 1687 22
rect 1683 18 1687 20
rect 1692 22 1698 23
rect 1692 20 1694 22
rect 1696 20 1698 22
rect 1692 13 1698 20
rect 1722 22 1726 24
rect 1722 20 1723 22
rect 1725 20 1726 22
rect 1722 15 1726 20
rect 1730 22 1734 33
rect 1738 36 1754 39
rect 1738 34 1739 36
rect 1741 35 1754 36
rect 1741 34 1742 35
rect 1738 29 1742 34
rect 1862 63 1868 69
rect 1823 62 1843 63
rect 1823 60 1839 62
rect 1841 60 1843 62
rect 1862 61 1864 63
rect 1866 61 1868 63
rect 1862 60 1868 61
rect 1875 60 1879 62
rect 1823 59 1843 60
rect 1738 27 1739 29
rect 1741 27 1742 29
rect 1738 25 1742 27
rect 1775 55 1793 56
rect 1775 53 1789 55
rect 1791 53 1793 55
rect 1775 52 1793 53
rect 1775 46 1779 52
rect 1811 56 1812 58
rect 1823 55 1827 59
rect 1875 58 1876 60
rect 1878 58 1879 60
rect 1775 44 1776 46
rect 1778 44 1779 46
rect 1771 23 1772 34
rect 1775 31 1779 44
rect 1794 39 1800 40
rect 1775 27 1790 31
rect 1786 23 1790 27
rect 1815 51 1827 55
rect 1815 46 1819 51
rect 1815 44 1816 46
rect 1818 44 1819 46
rect 1815 32 1819 44
rect 1849 55 1853 57
rect 1849 53 1850 55
rect 1852 53 1853 55
rect 1849 47 1853 53
rect 1875 55 1879 58
rect 1875 51 1899 55
rect 1849 43 1860 47
rect 1856 37 1860 43
rect 1895 47 1899 51
rect 1875 46 1891 47
rect 1875 44 1887 46
rect 1889 44 1891 46
rect 1875 43 1891 44
rect 1895 45 1900 47
rect 1895 43 1897 45
rect 1899 43 1900 45
rect 1875 37 1879 43
rect 1895 41 1900 43
rect 1895 39 1899 41
rect 1856 36 1879 37
rect 1856 34 1858 36
rect 1860 34 1879 36
rect 1856 33 1879 34
rect 1815 29 1832 32
rect 1815 28 1829 29
rect 1828 27 1829 28
rect 1831 27 1832 29
rect 1817 24 1823 25
rect 1730 21 1763 22
rect 1730 19 1759 21
rect 1761 19 1763 21
rect 1730 18 1763 19
rect 1786 22 1803 23
rect 1786 20 1799 22
rect 1801 20 1803 22
rect 1786 19 1803 20
rect 1817 22 1819 24
rect 1821 22 1823 24
rect 1722 13 1723 15
rect 1725 13 1726 15
rect 1778 15 1784 16
rect 1778 13 1780 15
rect 1782 13 1784 15
rect 1817 13 1823 22
rect 1828 22 1832 27
rect 1828 20 1829 22
rect 1831 20 1832 22
rect 1828 18 1832 20
rect 1837 22 1843 23
rect 1837 20 1839 22
rect 1841 20 1843 22
rect 1837 13 1843 20
rect 1867 22 1871 24
rect 1867 20 1868 22
rect 1870 20 1871 22
rect 1867 15 1871 20
rect 1875 22 1879 33
rect 1883 36 1899 39
rect 1883 34 1884 36
rect 1886 35 1899 36
rect 1886 34 1887 35
rect 1883 29 1887 34
rect 1883 27 1884 29
rect 1886 27 1887 29
rect 1883 25 1887 27
rect 1967 63 1973 69
rect 1928 62 1948 63
rect 1928 60 1944 62
rect 1946 60 1948 62
rect 1967 61 1969 63
rect 1971 61 1973 63
rect 1967 60 1973 61
rect 1980 60 1984 62
rect 1928 59 1948 60
rect 1916 56 1917 58
rect 1928 55 1932 59
rect 1980 58 1981 60
rect 1983 58 1984 60
rect 1920 51 1932 55
rect 1920 46 1924 51
rect 1920 44 1921 46
rect 1923 44 1924 46
rect 1920 32 1924 44
rect 1954 55 1958 57
rect 1954 53 1955 55
rect 1957 53 1958 55
rect 1954 47 1958 53
rect 1980 55 1984 58
rect 1980 51 2004 55
rect 1954 43 1965 47
rect 1961 37 1965 43
rect 2000 47 2004 51
rect 1980 46 1996 47
rect 1980 44 1992 46
rect 1994 44 1996 46
rect 1980 43 1996 44
rect 2000 45 2005 47
rect 2000 43 2002 45
rect 2004 43 2005 45
rect 1980 37 1984 43
rect 2000 41 2005 43
rect 2000 39 2004 41
rect 1961 36 1984 37
rect 1961 34 1963 36
rect 1965 34 1984 36
rect 1961 33 1984 34
rect 1920 29 1937 32
rect 1920 28 1934 29
rect 1933 27 1934 28
rect 1936 27 1937 29
rect 1922 24 1928 25
rect 1922 22 1924 24
rect 1926 22 1928 24
rect 1875 21 1908 22
rect 1875 19 1904 21
rect 1906 19 1908 21
rect 1875 18 1908 19
rect 1867 13 1868 15
rect 1870 13 1871 15
rect 1922 13 1928 22
rect 1933 22 1937 27
rect 1933 20 1934 22
rect 1936 20 1937 22
rect 1933 18 1937 20
rect 1942 22 1948 23
rect 1942 20 1944 22
rect 1946 20 1948 22
rect 1942 13 1948 20
rect 1972 22 1976 24
rect 1972 20 1973 22
rect 1975 20 1976 22
rect 1972 15 1976 20
rect 1980 22 1984 33
rect 1988 36 2004 39
rect 1988 34 1989 36
rect 1991 35 2004 36
rect 1991 34 1992 35
rect 1988 29 1992 34
rect 1988 27 1989 29
rect 1991 27 1992 29
rect 1988 25 1992 27
rect 1980 21 2013 22
rect 1980 19 2009 21
rect 2011 19 2013 21
rect 1980 18 2013 19
rect 1972 13 1973 15
rect 1975 13 1976 15
<< via1 >>
rect 51 198 53 200
rect 66 207 68 209
rect 91 198 93 200
rect 34 182 36 184
rect 74 183 76 185
rect 105 184 107 186
rect 167 207 169 209
rect 121 192 123 194
rect 194 207 196 209
rect 218 195 220 197
rect 186 184 188 186
rect 365 187 367 189
rect 379 197 381 199
rect 421 197 423 199
rect 396 180 398 182
rect 404 189 406 191
rect 436 206 438 208
rect 444 198 446 200
rect 468 206 470 208
rect 495 206 497 208
rect 492 173 494 175
rect 570 184 572 186
rect 584 197 586 199
rect 626 197 628 199
rect 601 180 603 182
rect 609 189 611 191
rect 641 206 643 208
rect 649 196 651 198
rect 673 206 675 208
rect 700 206 702 208
rect 697 173 699 175
rect 1841 198 1843 200
rect 746 180 748 182
rect 1856 207 1858 209
rect 1881 198 1883 200
rect 1824 182 1826 184
rect 1864 183 1866 185
rect 1895 184 1897 186
rect 1957 207 1959 209
rect 1984 207 1986 209
rect 2008 195 2010 197
rect 1976 184 1978 186
rect 66 135 68 137
rect 35 119 37 121
rect 74 126 76 128
rect 49 118 51 120
rect 91 118 93 120
rect 106 109 108 111
rect 162 142 164 144
rect 114 117 116 119
rect 138 109 140 111
rect 165 109 167 111
rect 211 108 213 110
rect 238 107 240 109
rect 262 109 264 111
rect 289 109 291 111
rect 364 133 366 135
rect 381 117 383 119
rect 404 132 406 134
rect 396 108 398 110
rect 421 117 423 119
rect 435 131 437 133
rect 335 102 337 104
rect 516 131 518 133
rect 497 108 499 110
rect 524 108 526 110
rect 569 133 571 135
rect 548 120 550 122
rect 586 117 588 119
rect 609 132 611 134
rect 601 108 603 110
rect 626 117 628 119
rect 640 131 642 133
rect 721 131 723 133
rect 656 116 658 118
rect 702 108 704 110
rect 729 108 731 110
rect 753 120 755 122
rect 808 135 810 137
rect 858 126 860 128
rect 840 109 842 111
rect 867 109 869 111
rect 913 109 915 111
rect 922 135 924 137
rect 955 127 957 129
rect 945 109 947 111
rect 972 109 974 111
rect 1058 135 1060 137
rect 1026 127 1028 129
rect 1018 102 1020 104
rect 1090 109 1092 111
rect 1117 109 1119 111
rect 1163 109 1165 111
rect 1172 135 1174 137
rect 1207 127 1209 129
rect 1195 109 1197 111
rect 1222 109 1224 111
rect 1308 135 1310 137
rect 1276 127 1278 129
rect 1268 103 1270 105
rect 1340 109 1342 111
rect 1367 109 1369 111
rect 1413 109 1415 111
rect 1422 135 1424 137
rect 1457 127 1459 129
rect 1445 109 1447 111
rect 1472 109 1474 111
rect 1558 135 1560 137
rect 1526 127 1528 129
rect 1518 103 1520 105
rect 1608 126 1610 128
rect 1590 109 1592 111
rect 1617 109 1619 111
rect 1663 109 1665 111
rect 1672 135 1674 137
rect 1695 109 1697 111
rect 1722 109 1724 111
rect 1768 102 1770 104
rect 1856 135 1858 137
rect 1864 126 1866 128
rect 1839 118 1841 120
rect 1881 118 1883 120
rect 1896 109 1898 111
rect 1952 142 1954 144
rect 1904 117 1906 119
rect 1928 109 1930 111
rect 1955 109 1957 111
rect 2001 106 2003 108
rect 939 71 941 73
rect 1110 71 1112 73
rect 1360 70 1362 72
rect 1949 71 1951 73
rect 40 27 42 29
rect 72 53 74 55
rect 99 53 101 55
rect 71 36 73 38
rect 145 53 147 55
rect 177 53 179 55
rect 154 27 156 29
rect 204 53 206 55
rect 187 35 189 37
rect 258 35 260 37
rect 290 27 292 29
rect 322 53 324 55
rect 349 53 351 55
rect 321 36 323 38
rect 395 53 397 55
rect 427 53 429 55
rect 404 27 406 29
rect 454 53 456 55
rect 439 35 441 37
rect 508 35 510 37
rect 540 27 542 29
rect 572 53 574 55
rect 599 53 601 55
rect 645 53 647 55
rect 597 19 599 21
rect 677 53 679 55
rect 654 27 656 29
rect 704 53 706 55
rect 689 35 691 37
rect 758 35 760 37
rect 790 27 792 29
rect 822 53 824 55
rect 849 53 851 55
rect 895 53 897 55
rect 856 43 858 45
rect 847 19 849 21
rect 927 53 929 55
rect 904 27 906 29
rect 954 53 956 55
rect 939 36 941 38
rect 1050 27 1052 29
rect 1082 53 1084 55
rect 1109 53 1111 55
rect 1094 35 1096 37
rect 1155 53 1157 55
rect 1245 60 1247 62
rect 1187 53 1189 55
rect 1164 27 1166 29
rect 1214 53 1216 55
rect 1197 35 1199 37
rect 1268 35 1270 37
rect 1300 27 1302 29
rect 1332 53 1334 55
rect 1359 53 1361 55
rect 1345 35 1347 37
rect 1405 53 1407 55
rect 1437 53 1439 55
rect 1414 27 1416 29
rect 1464 53 1466 55
rect 1449 35 1451 37
rect 1510 43 1512 45
rect 1518 35 1520 37
rect 1550 27 1552 29
rect 1582 53 1584 55
rect 1609 53 1611 55
rect 1582 36 1584 38
rect 1655 53 1657 55
rect 1687 53 1689 55
rect 1664 27 1666 29
rect 1714 53 1716 55
rect 1699 35 1701 37
rect 1768 35 1770 37
rect 1800 27 1802 29
rect 1832 53 1834 55
rect 1859 53 1861 55
rect 1832 36 1834 38
rect 1905 53 1907 55
rect 1937 53 1939 55
rect 1914 27 1916 29
rect 1964 53 1966 55
rect 1949 36 1951 38
<< via2 >>
rect 445 219 447 221
rect 35 114 37 116
rect 121 192 123 194
rect 121 176 123 178
rect 126 157 128 159
rect 365 202 367 204
rect 114 117 116 119
rect 444 198 446 200
rect 570 184 572 186
rect 860 206 862 208
rect 875 194 877 196
rect 874 168 876 170
rect 874 145 876 147
rect 858 126 860 128
rect 656 116 658 118
rect 874 121 876 123
rect 1018 117 1020 119
rect 35 89 37 91
rect 114 88 116 90
rect 221 89 223 91
rect 1608 126 1610 128
rect 1049 117 1051 119
rect 889 103 891 105
rect 256 89 258 91
rect 656 99 658 101
rect 1008 93 1010 95
rect 1032 93 1034 95
rect 1257 88 1259 90
rect 1282 88 1284 90
rect 1503 90 1505 92
rect 1904 117 1906 119
rect 1528 90 1530 92
rect 1904 100 1906 102
rect 1801 89 1803 91
rect 939 61 941 63
rect 1082 71 1084 73
rect 1101 61 1103 63
rect 1345 64 1347 66
rect 1121 61 1123 63
rect 939 45 941 47
rect 1801 73 1803 75
rect 1949 61 1951 63
rect 1949 45 1951 47
rect 1082 35 1084 37
rect 1345 35 1347 37
rect 597 19 599 21
<< labels >>
rlabel alu1 936 29 936 29 5 Vss
rlabel alu1 9 38 9 38 5 c2
rlabel alu1 98 21 98 21 5 p33
rlabel alu1 348 21 348 21 5 p32
rlabel alu1 598 21 598 21 5 p31
rlabel alu1 607 46 607 46 5 s13
rlabel alu1 848 21 848 21 5 p30
rlabel alu1 857 46 857 46 5 s12
rlabel alu1 1001 42 1001 42 5 r4
rlabel alu1 751 42 751 42 5 r5
rlabel alu1 501 42 501 42 5 r6
rlabel alu1 251 42 251 42 5 r7
rlabel alu1 357 46 357 46 5 sha
rlabel alu1 107 46 107 46 5 cha
rlabel alu1 1867 46 1867 46 5 p02
rlabel alu1 1858 21 1858 21 5 s00
rlabel alu1 1617 46 1617 46 5 p03
rlabel alu1 1608 21 1608 21 5 s01
rlabel alu1 1367 46 1367 46 5 Vss
rlabel alu1 1358 21 1358 21 5 s02
rlabel alu1 1117 46 1117 46 5 Vss
rlabel alu1 1108 21 1108 21 5 s03
rlabel alu1 1019 38 1019 38 5 c1
rlabel alu1 1261 42 1261 42 5 s13
rlabel alu1 1511 42 1511 42 5 s12
rlabel alu1 1946 29 1946 29 5 Vss
rlabel alu1 122 196 122 196 1 p31
rlabel alu1 212 122 212 122 1 p32
rlabel alu1 115 117 115 117 1 p33
rlabel alu1 35 119 35 119 1 p30
rlabel alu1 43 205 43 205 1 a2
rlabel via1 35 183 35 183 1 b3
rlabel alu1 83 203 83 203 1 a3
rlabel alu1 83 191 83 191 1 b2
rlabel alu1 83 114 83 114 1 a3
rlabel alu1 75 135 75 135 1 b3
rlabel via1 67 135 67 135 1 b2
rlabel alu1 59 113 59 113 1 a2
rlabel alu1 239 117 239 117 1 cha
rlabel alu1 288 143 288 143 1 c1
rlabel alu1 271 135 271 135 1 c1
rlabel alu1 297 118 297 118 1 c0
rlabel alu1 263 115 263 115 1 c0
rlabel alu1 336 122 336 122 1 sha
rlabel alu1 452 121 452 121 5 p21
rlabel alu1 413 114 413 114 5 a3
rlabel alu1 373 112 373 112 5 a2
rlabel alu1 413 203 413 203 5 a3
rlabel alu1 389 204 389 204 5 a2
rlabel alu1 405 182 405 182 5 b1
rlabel via1 397 182 397 182 5 b0
rlabel alu1 413 126 413 126 5 b0
rlabel via1 365 134 365 134 5 b1
rlabel via1 570 134 570 134 5 b3
rlabel alu1 618 126 618 126 5 b2
rlabel alu1 610 182 610 182 5 b3
rlabel via1 602 182 602 182 5 b2
rlabel alu1 542 195 542 195 5 p22
rlabel alu1 445 200 445 200 5 p23
rlabel alu1 365 198 365 198 5 p20
rlabel alu1 657 121 657 121 5 p11
rlabel alu1 747 195 747 195 5 p12
rlabel alu1 570 198 570 198 5 p10
rlabel alu1 650 200 650 200 5 p13
rlabel alu1 594 204 594 204 5 a0
rlabel alu1 618 203 618 203 5 a1
rlabel alu1 618 114 618 114 5 a1
rlabel alu1 578 112 578 112 5 a0
rlabel alu1 1849 113 1849 113 1 a0
rlabel alu1 1857 135 1857 135 1 b0
rlabel alu1 1865 135 1865 135 1 b1
rlabel alu1 1873 114 1873 114 1 a1
rlabel alu1 1873 191 1873 191 1 b0
rlabel alu1 1873 203 1873 203 1 a1
rlabel alu1 1833 205 1833 205 1 a0
rlabel via1 1825 183 1825 183 1 b1
rlabel alu1 1825 119 1825 119 1 r0
rlabel alu1 1912 196 1912 196 1 r1
rlabel alu1 2002 122 2002 122 1 p02
rlabel alu1 1905 117 1905 117 1 p03
rlabel alu1 866 143 866 143 1 p23
rlabel alu1 1116 143 1116 143 1 p22
rlabel alu1 1125 118 1125 118 1 p12
rlabel alu1 1366 143 1366 143 1 p21
rlabel alu1 1375 118 1375 118 1 p11
rlabel alu1 1616 143 1616 143 1 p20
rlabel alu1 1625 118 1625 118 1 p10
rlabel alu1 1704 135 1704 135 5 Vss
rlabel alu1 777 126 777 126 5 c0
rlabel alu1 1019 122 1019 122 5 s03
rlabel alu1 1269 122 1269 122 5 s02
rlabel alu1 1519 122 1519 122 5 s01
rlabel alu1 1769 122 1769 122 5 s00
rlabel alu1 2011 42 2011 42 1 r2
rlabel alu1 1761 42 1761 42 1 r3
rlabel alu1 875 118 875 118 1 p13
rlabel alu1 1488 155 1488 155 1 Vdd
rlabel alu1 1905 159 1905 159 1 Vdd
rlabel alu1 1455 90 1455 90 1 Vss
rlabel alu1 1288 72 1288 72 1 Vss
rlabel alu1 1466 8 1466 8 1 Vdd
rlabel alu1 1578 227 1578 227 1 Vss
<< end >>
