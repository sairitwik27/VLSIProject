magic
tech scmos
timestamp 1199203470
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 13 65 35 67
rect 43 66 45 70
rect 50 66 52 70
rect 13 57 15 65
rect 23 57 25 61
rect 33 57 35 65
rect 13 36 15 39
rect 9 34 17 36
rect 23 35 25 39
rect 9 32 11 34
rect 13 32 17 34
rect 9 30 17 32
rect 2 24 8 26
rect 2 22 4 24
rect 6 22 8 24
rect 2 20 8 22
rect 15 21 17 30
rect 22 33 28 35
rect 33 34 35 39
rect 43 35 45 38
rect 50 35 52 38
rect 22 31 24 33
rect 26 31 28 33
rect 22 29 28 31
rect 39 33 45 35
rect 49 33 55 35
rect 25 21 27 29
rect 39 26 41 33
rect 49 31 51 33
rect 53 31 55 33
rect 49 29 55 31
rect 49 26 51 29
rect 35 24 41 26
rect 45 24 51 26
rect 35 21 37 24
rect 45 21 47 24
rect 4 4 6 20
rect 56 16 62 18
rect 56 14 58 16
rect 60 14 62 16
rect 56 12 62 14
rect 15 8 17 12
rect 25 8 27 12
rect 35 4 37 12
rect 45 8 47 12
rect 56 4 58 12
rect 4 2 58 4
<< ndif >>
rect 10 18 15 21
rect 8 16 15 18
rect 8 14 10 16
rect 12 14 15 16
rect 8 12 15 14
rect 17 16 25 21
rect 17 14 20 16
rect 22 14 25 16
rect 17 12 25 14
rect 27 19 35 21
rect 27 17 30 19
rect 32 17 35 19
rect 27 12 35 17
rect 37 17 45 21
rect 37 15 40 17
rect 42 15 45 17
rect 37 12 45 15
rect 47 18 52 21
rect 47 16 54 18
rect 47 14 50 16
rect 52 14 54 16
rect 47 12 54 14
<< pdif >>
rect 38 57 43 66
rect 8 51 13 57
rect 6 49 13 51
rect 6 47 8 49
rect 10 47 13 49
rect 6 45 13 47
rect 8 39 13 45
rect 15 55 23 57
rect 15 53 18 55
rect 20 53 23 55
rect 15 48 23 53
rect 15 46 18 48
rect 20 46 23 48
rect 15 39 23 46
rect 25 50 33 57
rect 25 48 28 50
rect 30 48 33 50
rect 25 43 33 48
rect 25 41 28 43
rect 30 41 33 43
rect 25 39 33 41
rect 35 49 43 57
rect 35 47 38 49
rect 40 47 43 49
rect 35 39 43 47
rect 38 38 43 39
rect 45 38 50 66
rect 52 64 60 66
rect 52 62 55 64
rect 57 62 60 64
rect 52 57 60 62
rect 52 55 55 57
rect 57 55 60 57
rect 52 38 60 55
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 66 67
rect -2 64 66 65
rect 36 49 62 50
rect 36 47 38 49
rect 40 47 62 49
rect 36 46 62 47
rect 10 38 23 42
rect 10 34 14 38
rect 10 32 11 34
rect 13 32 14 34
rect 10 29 14 32
rect 18 33 31 34
rect 18 31 24 33
rect 26 31 31 33
rect 18 30 31 31
rect 18 21 22 30
rect 58 26 62 46
rect 41 22 62 26
rect 41 18 45 22
rect 38 17 45 18
rect 38 15 40 17
rect 42 15 45 17
rect 38 14 45 15
rect -2 0 66 8
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 15 12 17 21
rect 25 12 27 21
rect 35 12 37 21
rect 45 12 47 21
<< pmos >>
rect 13 39 15 57
rect 23 39 25 57
rect 33 39 35 57
rect 43 38 45 66
rect 50 38 52 66
<< polyct0 >>
rect 4 22 6 24
rect 51 31 53 33
rect 58 14 60 16
<< polyct1 >>
rect 11 32 13 34
rect 24 31 26 33
<< ndifct0 >>
rect 10 14 12 16
rect 20 14 22 16
rect 30 17 32 19
rect 50 14 52 16
<< ndifct1 >>
rect 40 15 42 17
<< ntiect1 >>
rect 5 65 7 67
<< pdifct0 >>
rect 8 47 10 49
rect 18 53 20 55
rect 18 46 20 48
rect 28 48 30 50
rect 28 41 30 43
rect 55 62 57 64
rect 55 55 57 57
<< pdifct1 >>
rect 38 47 40 49
<< alu0 >>
rect 16 55 22 64
rect 16 53 18 55
rect 20 53 22 55
rect 53 62 55 64
rect 57 62 59 64
rect 53 57 59 62
rect 53 55 55 57
rect 57 55 59 57
rect 53 54 59 55
rect 2 49 12 50
rect 2 47 8 49
rect 10 47 12 49
rect 2 46 12 47
rect 16 48 22 53
rect 16 46 18 48
rect 20 46 22 48
rect 2 26 6 46
rect 16 45 22 46
rect 27 50 31 52
rect 27 48 28 50
rect 30 48 31 50
rect 27 43 31 48
rect 27 41 28 43
rect 30 42 31 43
rect 30 41 38 42
rect 27 38 38 41
rect 34 34 38 38
rect 34 33 55 34
rect 34 31 51 33
rect 53 31 55 33
rect 34 30 55 31
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 34 26 38 30
rect 29 22 38 26
rect 29 19 33 22
rect 2 16 14 17
rect 2 14 10 16
rect 12 14 14 16
rect 2 13 14 14
rect 19 16 23 18
rect 19 14 20 16
rect 22 14 23 16
rect 29 17 30 19
rect 32 17 33 19
rect 29 15 33 17
rect 48 16 62 17
rect 48 14 50 16
rect 52 14 58 16
rect 60 14 62 16
rect 19 8 23 14
rect 48 13 62 14
<< labels >>
rlabel alu0 8 15 8 15 6 bn
rlabel alu0 7 48 7 48 6 bn
rlabel alu0 4 31 4 31 6 bn
rlabel alu0 31 20 31 20 6 an
rlabel alu0 29 45 29 45 6 an
rlabel alu0 55 15 55 15 6 bn
rlabel alu0 44 32 44 32 6 an
rlabel alu1 12 32 12 32 6 b
rlabel alu1 28 32 28 32 6 a
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 40 20 40 6 b
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 24 52 24 6 z
rlabel alu1 60 36 60 36 6 z
rlabel alu1 52 48 52 48 6 z
<< end >>
