magic
tech scmos
timestamp 1608973463
<< ab >>
rect 5 4 45 76
rect 47 4 110 76
<< nwell >>
rect 0 36 115 81
<< pwell >>
rect 0 -1 115 36
<< poly >>
rect 63 70 65 74
rect 14 61 16 65
rect 24 63 26 68
rect 34 63 36 68
rect 14 39 16 43
rect 24 39 26 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 48 45 54 47
rect 48 43 50 45
rect 52 43 54 45
rect 99 70 101 74
rect 79 61 81 65
rect 89 61 91 65
rect 48 41 54 43
rect 14 37 20 39
rect 14 35 16 37
rect 18 35 20 37
rect 14 33 20 35
rect 24 37 30 39
rect 24 35 26 37
rect 28 35 30 37
rect 24 33 30 35
rect 14 28 16 33
rect 27 28 29 33
rect 34 28 36 41
rect 52 40 54 41
rect 63 40 65 43
rect 79 40 81 43
rect 52 38 65 40
rect 71 38 81 40
rect 89 39 91 43
rect 99 40 101 43
rect 55 30 57 38
rect 71 34 73 38
rect 64 32 73 34
rect 85 37 91 39
rect 85 35 87 37
rect 89 35 91 37
rect 85 33 91 35
rect 95 38 101 40
rect 95 36 97 38
rect 99 36 101 38
rect 95 34 101 36
rect 64 30 66 32
rect 68 30 73 32
rect 14 15 16 19
rect 64 28 73 30
rect 89 30 91 33
rect 71 25 73 28
rect 81 25 83 29
rect 89 28 93 30
rect 91 25 93 28
rect 98 25 100 34
rect 55 18 57 21
rect 27 12 29 17
rect 34 12 36 17
rect 55 16 60 18
rect 58 8 60 16
rect 71 12 73 16
rect 81 8 83 16
rect 91 8 93 13
rect 98 8 100 13
rect 58 6 83 8
<< ndif >>
rect 48 28 55 30
rect 9 25 14 28
rect 7 23 14 25
rect 7 21 9 23
rect 11 21 14 23
rect 7 19 14 21
rect 16 19 27 28
rect 18 17 27 19
rect 29 17 34 28
rect 36 23 41 28
rect 48 26 50 28
rect 52 26 55 28
rect 48 24 55 26
rect 36 21 43 23
rect 50 21 55 24
rect 57 25 62 30
rect 57 21 71 25
rect 36 19 39 21
rect 41 19 43 21
rect 36 17 43 19
rect 62 20 71 21
rect 62 18 64 20
rect 66 18 71 20
rect 18 11 25 17
rect 62 16 71 18
rect 73 23 81 25
rect 73 21 76 23
rect 78 21 81 23
rect 73 16 81 21
rect 83 21 91 25
rect 83 19 86 21
rect 88 19 91 21
rect 83 16 91 19
rect 18 9 20 11
rect 22 9 25 11
rect 18 7 25 9
rect 86 13 91 16
rect 93 13 98 25
rect 100 13 108 25
rect 102 11 108 13
rect 102 9 104 11
rect 106 9 108 11
rect 102 7 108 9
<< pdif >>
rect 18 61 24 63
rect 9 56 14 61
rect 7 54 14 56
rect 7 52 9 54
rect 11 52 14 54
rect 7 47 14 52
rect 7 45 9 47
rect 11 45 14 47
rect 7 43 14 45
rect 16 59 24 61
rect 16 57 19 59
rect 21 57 24 59
rect 16 50 24 57
rect 26 61 34 63
rect 26 59 29 61
rect 31 59 34 61
rect 26 54 34 59
rect 26 52 29 54
rect 31 52 34 54
rect 26 50 34 52
rect 36 61 43 63
rect 36 59 39 61
rect 41 59 43 61
rect 36 50 43 59
rect 16 43 22 50
rect 58 49 63 70
rect 56 47 63 49
rect 56 45 58 47
rect 60 45 63 47
rect 56 43 63 45
rect 65 68 77 70
rect 65 66 68 68
rect 70 66 77 68
rect 65 61 77 66
rect 94 61 99 70
rect 65 59 68 61
rect 70 59 79 61
rect 65 43 79 59
rect 81 54 89 61
rect 81 52 84 54
rect 86 52 89 54
rect 81 47 89 52
rect 81 45 84 47
rect 86 45 89 47
rect 81 43 89 45
rect 91 54 99 61
rect 91 52 94 54
rect 96 52 99 54
rect 91 43 99 52
rect 101 64 106 70
rect 101 62 108 64
rect 101 60 104 62
rect 106 60 108 62
rect 101 58 108 60
rect 101 43 106 58
<< alu1 >>
rect 3 71 112 76
rect 3 69 10 71
rect 12 69 84 71
rect 86 69 112 71
rect 3 68 112 69
rect 7 54 12 56
rect 7 52 9 54
rect 11 52 12 54
rect 48 57 60 63
rect 7 47 12 52
rect 7 45 9 47
rect 11 45 12 47
rect 7 43 12 45
rect 7 23 11 43
rect 39 48 43 55
rect 48 48 53 57
rect 39 46 53 48
rect 30 45 53 46
rect 30 43 36 45
rect 38 43 50 45
rect 52 43 53 45
rect 30 42 43 43
rect 47 42 53 43
rect 48 41 53 42
rect 22 37 36 38
rect 22 35 26 37
rect 28 35 36 37
rect 22 34 36 35
rect 7 21 9 23
rect 11 21 19 23
rect 7 17 19 21
rect 31 28 36 34
rect 31 26 32 28
rect 34 26 36 28
rect 31 25 36 26
rect 64 32 69 39
rect 92 54 108 55
rect 92 52 94 54
rect 96 52 108 54
rect 92 50 108 52
rect 64 31 66 32
rect 56 30 66 31
rect 68 30 69 32
rect 56 28 69 30
rect 56 26 59 28
rect 61 26 69 28
rect 56 25 69 26
rect 104 22 108 50
rect 84 21 108 22
rect 84 19 86 21
rect 88 19 108 21
rect 84 18 108 19
rect 3 11 112 12
rect 3 9 10 11
rect 12 9 20 11
rect 22 9 51 11
rect 53 9 104 11
rect 106 9 112 11
rect 3 4 112 9
<< alu2 >>
rect 31 28 64 29
rect 31 26 32 28
rect 34 26 59 28
rect 61 26 64 28
rect 31 25 64 26
<< ptie >>
rect 8 11 14 13
rect 8 9 10 11
rect 12 9 14 11
rect 8 7 14 9
rect 49 11 55 13
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< ntie >>
rect 8 71 14 73
rect 8 69 10 71
rect 12 69 14 71
rect 82 71 88 73
rect 8 67 14 69
rect 82 69 84 71
rect 86 69 88 71
rect 82 67 88 69
<< nmos >>
rect 14 19 16 28
rect 27 17 29 28
rect 34 17 36 28
rect 55 21 57 30
rect 71 16 73 25
rect 81 16 83 25
rect 91 13 93 25
rect 98 13 100 25
<< pmos >>
rect 14 43 16 61
rect 24 50 26 63
rect 34 50 36 63
rect 63 43 65 70
rect 79 43 81 61
rect 89 43 91 61
rect 99 43 101 70
<< polyct0 >>
rect 16 35 18 37
rect 87 35 89 37
rect 97 36 99 38
<< polyct1 >>
rect 36 43 38 45
rect 50 43 52 45
rect 26 35 28 37
rect 66 30 68 32
<< ndifct0 >>
rect 50 26 52 28
rect 39 19 41 21
rect 64 18 66 20
rect 76 21 78 23
<< ndifct1 >>
rect 9 21 11 23
rect 86 19 88 21
rect 20 9 22 11
rect 104 9 106 11
<< ntiect1 >>
rect 10 69 12 71
rect 84 69 86 71
<< ptiect1 >>
rect 10 9 12 11
rect 51 9 53 11
<< pdifct0 >>
rect 19 57 21 59
rect 29 59 31 61
rect 29 52 31 54
rect 39 59 41 61
rect 58 45 60 47
rect 68 66 70 68
rect 68 59 70 61
rect 84 52 86 54
rect 84 45 86 47
rect 104 60 106 62
<< pdifct1 >>
rect 9 52 11 54
rect 9 45 11 47
rect 94 52 96 54
<< alu0 >>
rect 17 59 23 68
rect 17 57 19 59
rect 21 57 23 59
rect 17 56 23 57
rect 28 61 32 63
rect 28 59 29 61
rect 31 59 32 61
rect 28 54 32 59
rect 37 61 43 68
rect 67 66 68 68
rect 70 66 71 68
rect 37 59 39 61
rect 41 59 43 61
rect 37 58 43 59
rect 67 61 71 66
rect 67 59 68 61
rect 70 59 71 61
rect 67 57 71 59
rect 75 62 108 63
rect 75 60 104 62
rect 106 60 108 62
rect 75 59 108 60
rect 28 53 29 54
rect 15 52 29 53
rect 31 52 32 54
rect 15 49 32 52
rect 15 37 19 49
rect 75 48 79 59
rect 56 47 79 48
rect 56 45 58 47
rect 60 45 79 47
rect 56 44 79 45
rect 56 38 60 44
rect 15 35 16 37
rect 18 35 19 37
rect 15 30 19 35
rect 15 26 27 30
rect 11 23 12 25
rect 23 22 27 26
rect 49 34 60 38
rect 49 28 53 34
rect 75 38 79 44
rect 83 54 87 56
rect 83 52 84 54
rect 86 52 87 54
rect 83 47 87 52
rect 83 45 84 47
rect 86 46 87 47
rect 86 45 99 46
rect 83 42 99 45
rect 95 40 99 42
rect 95 38 100 40
rect 75 37 91 38
rect 75 35 87 37
rect 89 35 91 37
rect 75 34 91 35
rect 95 36 97 38
rect 99 36 100 38
rect 95 34 100 36
rect 49 26 50 28
rect 52 26 53 28
rect 49 24 53 26
rect 95 30 99 34
rect 75 26 99 30
rect 75 23 79 26
rect 23 21 43 22
rect 75 21 76 23
rect 78 21 79 23
rect 23 19 39 21
rect 41 19 43 21
rect 23 18 43 19
rect 62 20 68 21
rect 62 18 64 20
rect 66 18 68 20
rect 75 19 79 21
rect 62 12 68 18
<< via1 >>
rect 32 26 34 28
rect 59 26 61 28
<< labels >>
rlabel alu1 49 72 49 72 1 Vdd
rlabel alu1 25 72 25 72 6 vdd
rlabel alu1 47 7 47 7 1 Vss
rlabel alu1 106 39 106 39 1 sha
rlabel alu1 33 32 33 32 1 c0
rlabel alu1 67 35 67 35 1 c0
rlabel alu1 41 52 41 52 1 c1
rlabel alu1 58 60 58 60 1 c1
rlabel alu1 9 34 9 34 1 cha
<< end >>
