magic
tech scmos
timestamp 1608381361
<< ab >>
rect -36 5 4 77
rect 6 5 69 77
<< nwell >>
rect -41 37 74 82
<< pwell >>
rect -41 0 74 37
<< poly >>
rect 22 71 24 75
rect -27 62 -25 66
rect -17 64 -15 69
rect -7 64 -5 69
rect -27 40 -25 44
rect -17 40 -15 51
rect -7 48 -5 51
rect -7 46 -1 48
rect -7 44 -5 46
rect -3 44 -1 46
rect -7 42 -1 44
rect 7 46 13 48
rect 7 44 9 46
rect 11 44 13 46
rect 58 71 60 75
rect 38 62 40 66
rect 48 62 50 66
rect 7 42 13 44
rect -27 38 -21 40
rect -27 36 -25 38
rect -23 36 -21 38
rect -27 34 -21 36
rect -17 38 -11 40
rect -17 36 -15 38
rect -13 36 -11 38
rect -17 34 -11 36
rect -27 29 -25 34
rect -14 29 -12 34
rect -7 29 -5 42
rect 11 41 13 42
rect 22 41 24 44
rect 38 41 40 44
rect 11 39 24 41
rect 30 39 40 41
rect 48 40 50 44
rect 58 41 60 44
rect 14 31 16 39
rect 30 35 32 39
rect 23 33 32 35
rect 44 38 50 40
rect 44 36 46 38
rect 48 36 50 38
rect 44 34 50 36
rect 54 39 60 41
rect 54 37 56 39
rect 58 37 60 39
rect 54 35 60 37
rect 23 31 25 33
rect 27 31 32 33
rect -27 16 -25 20
rect 23 29 32 31
rect 48 31 50 34
rect 30 26 32 29
rect 40 26 42 30
rect 48 29 52 31
rect 50 26 52 29
rect 57 26 59 35
rect 14 19 16 22
rect -14 13 -12 18
rect -7 13 -5 18
rect 14 17 19 19
rect 17 9 19 17
rect 30 13 32 17
rect 40 9 42 17
rect 50 9 52 14
rect 57 9 59 14
rect 17 7 42 9
<< ndif >>
rect 7 29 14 31
rect -32 26 -27 29
rect -34 24 -27 26
rect -34 22 -32 24
rect -30 22 -27 24
rect -34 20 -27 22
rect -25 20 -14 29
rect -23 18 -14 20
rect -12 18 -7 29
rect -5 24 0 29
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect -5 22 2 24
rect 9 22 14 25
rect 16 26 21 31
rect 16 22 30 26
rect -5 20 -2 22
rect 0 20 2 22
rect -5 18 2 20
rect 21 21 30 22
rect 21 19 23 21
rect 25 19 30 21
rect -23 12 -16 18
rect 21 17 30 19
rect 32 24 40 26
rect 32 22 35 24
rect 37 22 40 24
rect 32 17 40 22
rect 42 22 50 26
rect 42 20 45 22
rect 47 20 50 22
rect 42 17 50 20
rect -23 10 -21 12
rect -19 10 -16 12
rect -23 8 -16 10
rect 45 14 50 17
rect 52 14 57 26
rect 59 14 67 26
rect 61 12 67 14
rect 61 10 63 12
rect 65 10 67 12
rect 61 8 67 10
<< pdif >>
rect -23 62 -17 64
rect -32 57 -27 62
rect -34 55 -27 57
rect -34 53 -32 55
rect -30 53 -27 55
rect -34 48 -27 53
rect -34 46 -32 48
rect -30 46 -27 48
rect -34 44 -27 46
rect -25 60 -17 62
rect -25 58 -22 60
rect -20 58 -17 60
rect -25 51 -17 58
rect -15 62 -7 64
rect -15 60 -12 62
rect -10 60 -7 62
rect -15 55 -7 60
rect -15 53 -12 55
rect -10 53 -7 55
rect -15 51 -7 53
rect -5 62 2 64
rect -5 60 -2 62
rect 0 60 2 62
rect -5 51 2 60
rect -25 44 -19 51
rect 17 50 22 71
rect 15 48 22 50
rect 15 46 17 48
rect 19 46 22 48
rect 15 44 22 46
rect 24 69 36 71
rect 24 67 27 69
rect 29 67 36 69
rect 24 62 36 67
rect 53 62 58 71
rect 24 60 27 62
rect 29 60 38 62
rect 24 44 38 60
rect 40 55 48 62
rect 40 53 43 55
rect 45 53 48 55
rect 40 48 48 53
rect 40 46 43 48
rect 45 46 48 48
rect 40 44 48 46
rect 50 55 58 62
rect 50 53 53 55
rect 55 53 58 55
rect 50 44 58 53
rect 60 65 65 71
rect 60 63 67 65
rect 60 61 63 63
rect 65 61 67 63
rect 60 59 67 61
rect 60 44 65 59
<< alu1 >>
rect -38 72 71 77
rect -38 70 -31 72
rect -29 70 43 72
rect 45 70 71 72
rect -38 69 71 70
rect -34 55 -29 57
rect -34 53 -32 55
rect -30 53 -29 55
rect 7 58 19 64
rect -34 48 -29 53
rect -34 46 -32 48
rect -30 46 -29 48
rect -34 44 -29 46
rect -34 24 -30 44
rect -2 49 2 56
rect 7 49 12 58
rect -2 47 12 49
rect -11 46 12 47
rect -11 44 -5 46
rect -3 44 9 46
rect 11 44 12 46
rect -11 43 2 44
rect 6 43 12 44
rect 7 42 12 43
rect -19 38 -5 39
rect -19 36 -15 38
rect -13 36 -5 38
rect -19 35 -5 36
rect -34 22 -32 24
rect -30 22 -22 24
rect -34 18 -22 22
rect -10 29 -5 35
rect -10 27 -9 29
rect -7 27 -5 29
rect -10 26 -5 27
rect 23 33 28 40
rect 51 55 67 56
rect 51 53 53 55
rect 55 53 67 55
rect 51 51 67 53
rect 23 32 25 33
rect 15 31 25 32
rect 27 31 28 33
rect 15 29 28 31
rect 15 27 18 29
rect 20 27 28 29
rect 15 26 28 27
rect 63 23 67 51
rect 43 22 67 23
rect 43 20 45 22
rect 47 20 67 22
rect 43 19 67 20
rect -38 12 71 13
rect -38 10 -31 12
rect -29 10 -21 12
rect -19 10 10 12
rect 12 10 63 12
rect 65 10 71 12
rect -38 5 71 10
<< alu2 >>
rect -10 29 23 30
rect -10 27 -9 29
rect -7 27 18 29
rect 20 27 23 29
rect -10 26 23 27
<< ptie >>
rect -33 12 -27 14
rect -33 10 -31 12
rect -29 10 -27 12
rect -33 8 -27 10
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
<< ntie >>
rect -33 72 -27 74
rect -33 70 -31 72
rect -29 70 -27 72
rect 41 72 47 74
rect -33 68 -27 70
rect 41 70 43 72
rect 45 70 47 72
rect 41 68 47 70
<< nmos >>
rect -27 20 -25 29
rect -14 18 -12 29
rect -7 18 -5 29
rect 14 22 16 31
rect 30 17 32 26
rect 40 17 42 26
rect 50 14 52 26
rect 57 14 59 26
<< pmos >>
rect -27 44 -25 62
rect -17 51 -15 64
rect -7 51 -5 64
rect 22 44 24 71
rect 38 44 40 62
rect 48 44 50 62
rect 58 44 60 71
<< polyct0 >>
rect -25 36 -23 38
rect 46 36 48 38
rect 56 37 58 39
<< polyct1 >>
rect -5 44 -3 46
rect 9 44 11 46
rect -15 36 -13 38
rect 25 31 27 33
<< ndifct0 >>
rect 9 27 11 29
rect -2 20 0 22
rect 23 19 25 21
rect 35 22 37 24
<< ndifct1 >>
rect -32 22 -30 24
rect 45 20 47 22
rect -21 10 -19 12
rect 63 10 65 12
<< ntiect1 >>
rect -31 70 -29 72
rect 43 70 45 72
<< ptiect1 >>
rect -31 10 -29 12
rect 10 10 12 12
<< pdifct0 >>
rect -22 58 -20 60
rect -12 60 -10 62
rect -12 53 -10 55
rect -2 60 0 62
rect 17 46 19 48
rect 27 67 29 69
rect 27 60 29 62
rect 43 53 45 55
rect 43 46 45 48
rect 63 61 65 63
<< pdifct1 >>
rect -32 53 -30 55
rect -32 46 -30 48
rect 53 53 55 55
<< alu0 >>
rect -24 60 -18 69
rect -24 58 -22 60
rect -20 58 -18 60
rect -24 57 -18 58
rect -13 62 -9 64
rect -13 60 -12 62
rect -10 60 -9 62
rect -13 55 -9 60
rect -4 62 2 69
rect 26 67 27 69
rect 29 67 30 69
rect -4 60 -2 62
rect 0 60 2 62
rect -4 59 2 60
rect 26 62 30 67
rect 26 60 27 62
rect 29 60 30 62
rect 26 58 30 60
rect 34 63 67 64
rect 34 61 63 63
rect 65 61 67 63
rect 34 60 67 61
rect -13 54 -12 55
rect -26 53 -12 54
rect -10 53 -9 55
rect -26 50 -9 53
rect -26 38 -22 50
rect 34 49 38 60
rect 15 48 38 49
rect 15 46 17 48
rect 19 46 38 48
rect 15 45 38 46
rect 15 39 19 45
rect -26 36 -25 38
rect -23 36 -22 38
rect -26 31 -22 36
rect -26 27 -14 31
rect -30 24 -29 26
rect -18 23 -14 27
rect 8 35 19 39
rect 8 29 12 35
rect 34 39 38 45
rect 42 55 46 57
rect 42 53 43 55
rect 45 53 46 55
rect 42 48 46 53
rect 42 46 43 48
rect 45 47 46 48
rect 45 46 58 47
rect 42 43 58 46
rect 54 41 58 43
rect 54 39 59 41
rect 34 38 50 39
rect 34 36 46 38
rect 48 36 50 38
rect 34 35 50 36
rect 54 37 56 39
rect 58 37 59 39
rect 54 35 59 37
rect 8 27 9 29
rect 11 27 12 29
rect 8 25 12 27
rect 54 31 58 35
rect 34 27 58 31
rect 34 24 38 27
rect -18 22 2 23
rect 34 22 35 24
rect 37 22 38 24
rect -18 20 -2 22
rect 0 20 2 22
rect -18 19 2 20
rect 21 21 27 22
rect 21 19 23 21
rect 25 19 27 21
rect 34 20 38 22
rect 21 13 27 19
<< via1 >>
rect -9 27 -7 29
rect 18 27 20 29
<< labels >>
rlabel alu1 17 61 17 61 6 b
rlabel alu1 8 73 8 73 1 Vdd
rlabel alu1 65 40 65 40 1 sum
rlabel alu1 -8 33 -8 33 6 a
rlabel alu1 -16 73 -16 73 6 vdd
rlabel alu1 0 53 0 53 6 b
rlabel alu1 6 8 6 8 1 Vss
rlabel alu1 26 36 26 36 1 a
rlabel alu1 -32 35 -32 35 1 cout
<< end >>
